* NGSPICE file created from wrapped_ibnalhaytham.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

.subckt wrapped_ibnalhaytham active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ user_clock2 vccd1 vssd1 wb_clk_i
XFILLER_28_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18869_ _18869_/A vssd1 vssd1 vccd1 vccd1 _26043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20900_ _20900_/A vssd1 vssd1 vccd1 vccd1 _20900_/X sky130_fd_sc_hd__clkbuf_1
X_21880_ _21912_/A vssd1 vssd1 vccd1 vccd1 _21880_/X sky130_fd_sc_hd__clkbuf_1
X_20831_ _20831_/A vssd1 vssd1 vccd1 vccd1 _20831_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20762_ _20754_/X _20755_/X _20756_/X _20757_/X _20758_/X _20759_/X vssd1 vssd1 vccd1
+ vccd1 _20763_/A sky130_fd_sc_hd__mux4_1
XFILLER_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23550_ _27764_/Q _27206_/Q _23559_/S vssd1 vssd1 vccd1 vccd1 _23551_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22501_ _22487_/X _22488_/X _22489_/X _22490_/X _22491_/X _22492_/X vssd1 vssd1 vccd1
+ vccd1 _22502_/A sky130_fd_sc_hd__mux4_1
XFILLER_39_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23481_ input24/X _23469_/X _23480_/X _23474_/X vssd1 vssd1 vccd1 vccd1 _27185_/D
+ sky130_fd_sc_hd__o211a_1
X_20693_ _20693_/A vssd1 vssd1 vccd1 vccd1 _20693_/X sky130_fd_sc_hd__clkbuf_1
X_22432_ _22432_/A vssd1 vssd1 vccd1 vccd1 _22432_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25220_ _25220_/A _25220_/B vssd1 vssd1 vccd1 vccd1 _25221_/B sky130_fd_sc_hd__xnor2_1
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22363_ _22347_/X _22348_/X _22349_/X _22350_/X _22352_/X _22354_/X vssd1 vssd1 vccd1
+ vccd1 _22364_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25151_ _25182_/A _25151_/B vssd1 vssd1 vccd1 vccd1 _25151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21314_ _21314_/A vssd1 vssd1 vccd1 vccd1 _21314_/X sky130_fd_sc_hd__clkbuf_1
X_24102_ _27399_/Q _24106_/B vssd1 vssd1 vccd1 vccd1 _24103_/A sky130_fd_sc_hd__and2_1
X_25082_ _25080_/X _25081_/X _25103_/S vssd1 vssd1 vccd1 vccd1 _25082_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22294_ _22294_/A vssd1 vssd1 vccd1 vccd1 _22294_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24033_ _24031_/X _24032_/X _24033_/S vssd1 vssd1 vccd1 vccd1 _24033_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21245_ _21231_/X _21234_/X _21237_/X _21240_/X _21241_/X _21242_/X vssd1 vssd1 vccd1
+ vccd1 _21246_/A sky130_fd_sc_hd__mux4_1
XFILLER_172_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21176_ _21176_/A vssd1 vssd1 vccd1 vccd1 _21176_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20127_ _20127_/A vssd1 vssd1 vccd1 vccd1 _20127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25984_ _25984_/CLK _25984_/D vssd1 vssd1 vccd1 vccd1 _25984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27723_ _27744_/CLK _27723_/D vssd1 vssd1 vccd1 vccd1 _27723_/Q sky130_fd_sc_hd__dfxtp_1
X_20058_ _20044_/X _20045_/X _20046_/X _20047_/X _20048_/X _20049_/X vssd1 vssd1 vccd1
+ vccd1 _20059_/A sky130_fd_sc_hd__mux4_1
X_24935_ _24935_/A vssd1 vssd1 vccd1 vccd1 _24935_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27654_ _27654_/CLK _27654_/D vssd1 vssd1 vccd1 vccd1 _27654_/Q sky130_fd_sc_hd__dfxtp_1
X_24866_ _24935_/A vssd1 vssd1 vccd1 vccd1 _24889_/A sky130_fd_sc_hd__clkbuf_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater190 _26012_/CLK vssd1 vssd1 vccd1 vccd1 _26013_/CLK sky130_fd_sc_hd__clkbuf_1
X_26605_ _21434_/X _26605_/D vssd1 vssd1 vccd1 vccd1 _26605_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_213 _14518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23817_ _23800_/X _23811_/X _23815_/X _23816_/X vssd1 vssd1 vccd1 vccd1 _27276_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 _14807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27585_ _27585_/CLK _27585_/D vssd1 vssd1 vccd1 vccd1 _27585_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24797_ _27632_/Q _24785_/X _24796_/Y _24787_/X vssd1 vssd1 vccd1 vccd1 _27632_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _17321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _27764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _26816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _15710_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14550_/Y sky130_fd_sc_hd__nor2_1
X_26536_ _21188_/X _26536_/D vssd1 vssd1 vccd1 vccd1 _26536_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_268 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23748_ _27786_/Q vssd1 vssd1 vccd1 vccd1 _23929_/A sky130_fd_sc_hd__buf_2
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_279 input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _27352_/Q _13450_/X _13451_/X _27320_/Q _13136_/X vssd1 vssd1 vccd1 vccd1
+ _14471_/A sky130_fd_sc_hd__a221oi_4
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14481_ _26633_/Q _14478_/X _14474_/X _14480_/Y vssd1 vssd1 vccd1 vccd1 _26633_/D
+ sky130_fd_sc_hd__a31o_1
X_26467_ _20948_/X _26467_/D vssd1 vssd1 vccd1 vccd1 _26467_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23679_ _24877_/A _27245_/Q _23683_/S vssd1 vssd1 vccd1 vccd1 _23680_/A sky130_fd_sc_hd__mux2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16220_ _16180_/X _16215_/X _16217_/Y _16218_/X _16219_/X vssd1 vssd1 vccd1 vccd1
+ _16357_/A sky130_fd_sc_hd__o41a_1
X_13432_ _13456_/A vssd1 vssd1 vccd1 vccd1 _13442_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25418_ _27747_/Q input59/X _25424_/S vssd1 vssd1 vccd1 vccd1 _25419_/A sky130_fd_sc_hd__mux2_1
X_26398_ _20699_/X _26398_/D vssd1 vssd1 vccd1 vccd1 _26398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _16151_/A _24301_/A vssd1 vssd1 vccd1 vccd1 _16301_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25349_ _25339_/B _25342_/A _25341_/Y _25339_/A vssd1 vssd1 vccd1 vccd1 _25350_/B
+ sky130_fd_sc_hd__o211a_1
X_13363_ _14753_/A vssd1 vssd1 vccd1 vccd1 _13363_/X sky130_fd_sc_hd__buf_2
XFILLER_127_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15102_ _15102_/A vssd1 vssd1 vccd1 vccd1 _26401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16082_ _16646_/B vssd1 vssd1 vccd1 vccd1 _16625_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13294_ _27013_/Q _13172_/X _13302_/S vssd1 vssd1 vccd1 vccd1 _13295_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15033_ _26431_/Q _15028_/X _15029_/X _15032_/Y vssd1 vssd1 vccd1 vccd1 _26431_/D
+ sky130_fd_sc_hd__a31o_1
X_27019_ _22868_/X _27019_/D vssd1 vssd1 vccd1 vccd1 _27019_/Q sky130_fd_sc_hd__dfxtp_1
X_19910_ _19898_/X _19899_/X _19900_/X _19901_/X _19903_/X _19905_/X vssd1 vssd1 vccd1
+ vccd1 _19911_/A sky130_fd_sc_hd__mux4_1
XFILLER_142_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19841_ _19841_/A vssd1 vssd1 vccd1 vccd1 _19841_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16984_ input37/X vssd1 vssd1 vccd1 vccd1 _17220_/A sky130_fd_sc_hd__buf_2
XFILLER_150_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19772_ _19764_/X _19765_/X _19766_/X _19767_/X _19768_/X _19769_/X vssd1 vssd1 vccd1
+ vccd1 _19773_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18723_ _18723_/A vssd1 vssd1 vccd1 vccd1 _26023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15935_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15935_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18654_ _18676_/A vssd1 vssd1 vccd1 vccd1 _18663_/S sky130_fd_sc_hd__buf_2
XFILLER_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15866_ _15868_/A vssd1 vssd1 vccd1 vccd1 _15866_/Y sky130_fd_sc_hd__inv_2
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17605_ _17605_/A vssd1 vssd1 vccd1 vccd1 _25875_/D sky130_fd_sc_hd__clkbuf_1
X_14817_ _14817_/A vssd1 vssd1 vccd1 vccd1 _26521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18585_ _27859_/Q _27194_/Q input5/X vssd1 vssd1 vccd1 vccd1 _18601_/A sky130_fd_sc_hd__or3_1
XFILLER_188_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15797_ _13086_/X _26100_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15798_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17536_ _17431_/X _25845_/Q _17540_/S vssd1 vssd1 vccd1 vccd1 _17537_/A sky130_fd_sc_hd__mux2_1
X_14748_ _14747_/X _26542_/Q _14757_/S vssd1 vssd1 vccd1 vccd1 _14749_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17467_ _17466_/X _25824_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17468_/A sky130_fd_sc_hd__mux2_1
X_14679_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14679_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19206_ _26697_/Q _26665_/Q _26633_/Q _26601_/Q _19179_/X _19087_/X vssd1 vssd1 vccd1
+ vccd1 _19206_/X sky130_fd_sc_hd__mux4_2
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16418_ _16708_/A _16708_/B vssd1 vssd1 vccd1 vccd1 _16732_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17398_ input73/X vssd1 vssd1 vccd1 vccd1 _20800_/A sky130_fd_sc_hd__inv_2
Xrepeater82 _27295_/CLK vssd1 vssd1 vccd1 vccd1 _27427_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_158_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater93 _25935_/CLK vssd1 vssd1 vccd1 vccd1 _26001_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_118_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19137_ _26822_/Q _26790_/Q _26758_/Q _26726_/Q _18913_/X _18930_/X vssd1 vssd1 vccd1
+ vccd1 _19137_/X sky130_fd_sc_hd__mux4_2
XFILLER_146_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16349_ _16753_/B _16349_/B vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__and2_1
XFILLER_173_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19068_ _24403_/A _19067_/X _24405_/A vssd1 vssd1 vccd1 vccd1 _19068_/X sky130_fd_sc_hd__o21a_1
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_528 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18019_ _18019_/A _17935_/X vssd1 vssd1 vccd1 vccd1 _18019_/X sky130_fd_sc_hd__or2b_1
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21030_ _21030_/A vssd1 vssd1 vccd1 vccd1 _21030_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22981_ _23029_/A vssd1 vssd1 vccd1 vccd1 _22981_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24720_ _27604_/Q _24714_/X _24719_/X _24717_/X vssd1 vssd1 vccd1 vccd1 _27604_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21932_ _21998_/A vssd1 vssd1 vccd1 vccd1 _21932_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24651_ _27578_/Q _24643_/X _24646_/X _24650_/X vssd1 vssd1 vccd1 vccd1 _27578_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21863_ _21911_/A vssd1 vssd1 vccd1 vccd1 _21863_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23602_ _23617_/A _23602_/B vssd1 vssd1 vccd1 vccd1 _23603_/A sky130_fd_sc_hd__and2_1
X_20814_ _20791_/X _20795_/X _20799_/X _20803_/X _20804_/X _20805_/X vssd1 vssd1 vccd1
+ vccd1 _20815_/A sky130_fd_sc_hd__mux4_1
X_27370_ _27372_/CLK _27370_/D vssd1 vssd1 vccd1 vccd1 _27370_/Q sky130_fd_sc_hd__dfxtp_1
X_21794_ _21826_/A vssd1 vssd1 vccd1 vccd1 _21794_/X sky130_fd_sc_hd__clkbuf_1
X_24582_ _24582_/A vssd1 vssd1 vccd1 vccd1 _27551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26321_ _20437_/X _26321_/D vssd1 vssd1 vccd1 vccd1 _26321_/Q sky130_fd_sc_hd__dfxtp_1
X_23533_ _24848_/A _27201_/Q _23542_/S vssd1 vssd1 vccd1 vccd1 _23534_/B sky130_fd_sc_hd__mux2_1
X_20745_ _20745_/A vssd1 vssd1 vccd1 vccd1 _20745_/X sky130_fd_sc_hd__clkbuf_1
X_26252_ _20195_/X _26252_/D vssd1 vssd1 vccd1 vccd1 _26252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23464_ input16/X _23455_/X _23463_/X _23461_/X vssd1 vssd1 vccd1 vccd1 _27178_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20676_ _20668_/X _20669_/X _20670_/X _20671_/X _20672_/X _20673_/X vssd1 vssd1 vccd1
+ vccd1 _20677_/A sky130_fd_sc_hd__mux4_1
XFILLER_137_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25203_ _25203_/A _25203_/B vssd1 vssd1 vccd1 vccd1 _25205_/A sky130_fd_sc_hd__nand2_1
XFILLER_195_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22415_ _22401_/X _22402_/X _22403_/X _22404_/X _22405_/X _22406_/X vssd1 vssd1 vccd1
+ vccd1 _22416_/A sky130_fd_sc_hd__mux4_1
XFILLER_52_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26183_ _19953_/X _26183_/D vssd1 vssd1 vccd1 vccd1 _26183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23395_ _27784_/Q _27264_/Q vssd1 vssd1 vccd1 vccd1 _23395_/X sky130_fd_sc_hd__xor2_1
XFILLER_52_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25134_ _27523_/Q _27491_/Q vssd1 vssd1 vccd1 vccd1 _25136_/A sky130_fd_sc_hd__and2_1
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22346_ _22346_/A vssd1 vssd1 vccd1 vccd1 _22346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22277_ _22261_/X _22262_/X _22263_/X _22264_/X _22266_/X _22268_/X vssd1 vssd1 vccd1
+ vccd1 _22278_/A sky130_fd_sc_hd__mux4_1
X_25065_ _27076_/Q _27108_/Q _25088_/S vssd1 vssd1 vccd1 vccd1 _25065_/X sky130_fd_sc_hd__mux2_1
X_24016_ _25939_/Q _26005_/Q _25838_/Q _26037_/Q _23993_/X _23976_/X vssd1 vssd1 vccd1
+ vccd1 _24016_/X sky130_fd_sc_hd__mux4_1
X_21228_ _21228_/A vssd1 vssd1 vccd1 vccd1 _21228_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21159_ _21144_/X _21146_/X _21148_/X _21150_/X _21151_/X _21152_/X vssd1 vssd1 vccd1
+ vccd1 _21160_/A sky130_fd_sc_hd__mux4_1
XFILLER_120_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13981_ _14356_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13981_/Y sky130_fd_sc_hd__nor2_1
X_25967_ _27326_/CLK _25967_/D vssd1 vssd1 vccd1 vccd1 _25967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15720_ _25075_/A vssd1 vssd1 vccd1 vccd1 _24980_/S sky130_fd_sc_hd__clkbuf_4
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27706_ _27706_/CLK _27706_/D vssd1 vssd1 vccd1 vccd1 _27706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_512 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24918_ _27773_/Q _24918_/B vssd1 vssd1 vccd1 vccd1 _24919_/B sky130_fd_sc_hd__nor2_1
X_12932_ _12932_/A vssd1 vssd1 vccd1 vccd1 _27859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25898_ _27153_/CLK _25898_/D vssd1 vssd1 vccd1 vccd1 _25898_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27637_ _27711_/CLK _27637_/D vssd1 vssd1 vccd1 vccd1 _27637_/Q sky130_fd_sc_hd__dfxtp_1
X_15651_ _15651_/A vssd1 vssd1 vccd1 vccd1 _26158_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24849_ _24863_/A _24849_/B vssd1 vssd1 vccd1 vccd1 _24849_/Y sky130_fd_sc_hd__nand2_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14602_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18370_ _26287_/Q _26255_/Q _26223_/Q _26191_/Q _17801_/X _17805_/X vssd1 vssd1 vccd1
+ vccd1 _18370_/X sky130_fd_sc_hd__mux4_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15582_ _26188_/Q _14753_/A _15584_/S vssd1 vssd1 vccd1 vccd1 _15583_/A sky130_fd_sc_hd__mux2_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27568_ _27568_/CLK _27568_/D vssd1 vssd1 vccd1 vccd1 _27568_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17319_/X _17320_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17321_/X sky130_fd_sc_hd__mux2_2
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _26618_/Q _14530_/X _14426_/B _14532_/Y vssd1 vssd1 vccd1 vccd1 _26618_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26519_ _21124_/X _26519_/D vssd1 vssd1 vccd1 vccd1 _26519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27499_ _27747_/CLK _27499_/D vssd1 vssd1 vccd1 vccd1 _27499_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _17252_/A vssd1 vssd1 vccd1 vccd1 _17252_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14464_ _14464_/A vssd1 vssd1 vccd1 vccd1 _15732_/A sky130_fd_sc_hd__buf_2
X_16203_ _27383_/Q vssd1 vssd1 vccd1 vccd1 _23035_/A sky130_fd_sc_hd__inv_2
XFILLER_168_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ _26972_/Q _13414_/X _13415_/S vssd1 vssd1 vccd1 vccd1 _13416_/A sky130_fd_sc_hd__mux2_1
X_17183_ _17181_/X _17182_/X _17159_/X vssd1 vssd1 vccd1 vccd1 _17183_/X sky130_fd_sc_hd__a21bo_1
X_14395_ _26658_/Q _14392_/X _14385_/X _14394_/Y vssd1 vssd1 vccd1 vccd1 _26658_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_155_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _16134_/A _16264_/B _16274_/C vssd1 vssd1 vccd1 vccd1 _16134_/X sky130_fd_sc_hd__or3_1
X_13346_ _13346_/A vssd1 vssd1 vccd1 vccd1 _26994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16065_ _16400_/A vssd1 vssd1 vccd1 vccd1 _16536_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_154_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ _13277_/A vssd1 vssd1 vccd1 vccd1 _27021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15016_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15016_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19824_ _19812_/X _19813_/X _19814_/X _19815_/X _19817_/X _19819_/X vssd1 vssd1 vccd1
+ vccd1 _19825_/A sky130_fd_sc_hd__mux4_1
XFILLER_190_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19755_ _19755_/A vssd1 vssd1 vccd1 vccd1 _19755_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16967_ _19313_/A _16967_/B _16967_/C vssd1 vssd1 vccd1 vccd1 _25907_/D sky130_fd_sc_hd__nand3_1
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18706_ _18706_/A vssd1 vssd1 vccd1 vccd1 _26015_/D sky130_fd_sc_hd__clkbuf_1
X_15918_ _15918_/A vssd1 vssd1 vccd1 vccd1 _15918_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16898_ _16309_/Y _16902_/A _16600_/Y _16093_/X vssd1 vssd1 vccd1 vccd1 _16898_/Y
+ sky130_fd_sc_hd__o31ai_1
X_19686_ _19678_/X _19679_/X _19680_/X _19681_/X _19682_/X _19683_/X vssd1 vssd1 vccd1
+ vccd1 _19687_/A sky130_fd_sc_hd__mux4_1
XFILLER_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15849_ _13228_/X _26076_/Q _15849_/S vssd1 vssd1 vccd1 vccd1 _15850_/A sky130_fd_sc_hd__mux2_1
X_18637_ _25985_/Q _17699_/X _18641_/S vssd1 vssd1 vccd1 vccd1 _18638_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18568_ _18566_/X _18567_/X _18568_/S vssd1 vssd1 vccd1 vccd1 _18568_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17519_ _17519_/A vssd1 vssd1 vccd1 vccd1 _25840_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18499_ _18379_/X _18496_/X _18498_/X _18384_/X vssd1 vssd1 vccd1 vccd1 _18499_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20530_ _20702_/A vssd1 vssd1 vccd1 vccd1 _20598_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20461_ _20461_/A vssd1 vssd1 vccd1 vccd1 _20461_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22200_ _22264_/A vssd1 vssd1 vccd1 vccd1 _22200_/X sky130_fd_sc_hd__clkbuf_1
X_23180_ _27129_/Q _17775_/X _23180_/S vssd1 vssd1 vccd1 vccd1 _23181_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20392_ _20424_/A vssd1 vssd1 vccd1 vccd1 _20392_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22131_ _22125_/X _22126_/X _22127_/X _22128_/X _22129_/X _22130_/X vssd1 vssd1 vccd1
+ vccd1 _22132_/A sky130_fd_sc_hd__mux4_1
XFILLER_145_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22062_ _22062_/A vssd1 vssd1 vccd1 vccd1 _22062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21013_ _21007_/X _21008_/X _21009_/X _21010_/X _21011_/X _21012_/X vssd1 vssd1 vccd1
+ vccd1 _21014_/A sky130_fd_sc_hd__mux4_1
XFILLER_88_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26870_ _22356_/X _26870_/D vssd1 vssd1 vccd1 vccd1 _26870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25821_ _26020_/CLK _25821_/D vssd1 vssd1 vccd1 vccd1 _25821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25752_ _25752_/A vssd1 vssd1 vccd1 vccd1 _27832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22964_ _22964_/A vssd1 vssd1 vccd1 vccd1 _22964_/X sky130_fd_sc_hd__clkbuf_1
X_24703_ _24729_/A vssd1 vssd1 vccd1 vccd1 _24703_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21915_ _22087_/A vssd1 vssd1 vccd1 vccd1 _21985_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25683_ _25673_/X _25674_/X _25675_/X _25676_/X _25677_/X _25678_/X vssd1 vssd1 vccd1
+ vccd1 _25684_/A sky130_fd_sc_hd__mux4_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22895_ _22943_/A vssd1 vssd1 vccd1 vccd1 _22895_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27422_ _27422_/CLK _27422_/D vssd1 vssd1 vccd1 vccd1 _27422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24634_ _24634_/A vssd1 vssd1 vccd1 vccd1 _27575_/D sky130_fd_sc_hd__clkbuf_1
X_21846_ _21912_/A vssd1 vssd1 vccd1 vccd1 _21846_/X sky130_fd_sc_hd__clkbuf_1
X_27353_ _27353_/CLK _27353_/D vssd1 vssd1 vccd1 vccd1 _27353_/Q sky130_fd_sc_hd__dfxtp_2
X_24565_ _27644_/Q _24565_/B vssd1 vssd1 vccd1 vccd1 _24566_/A sky130_fd_sc_hd__and2_1
X_21777_ _21825_/A vssd1 vssd1 vccd1 vccd1 _21777_/X sky130_fd_sc_hd__clkbuf_1
X_26304_ _20375_/X _26304_/D vssd1 vssd1 vccd1 vccd1 _26304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23516_ _27755_/Q vssd1 vssd1 vccd1 vccd1 _24831_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27284_ _27285_/CLK _27284_/D vssd1 vssd1 vccd1 vccd1 _27284_/Q sky130_fd_sc_hd__dfxtp_1
X_20728_ _20722_/X _20723_/X _20724_/X _20725_/X _20726_/X _20727_/X vssd1 vssd1 vccd1
+ vccd1 _20729_/A sky130_fd_sc_hd__mux4_1
XFILLER_12_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24496_ _24496_/A vssd1 vssd1 vccd1 vccd1 _27519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26235_ _20137_/X _26235_/D vssd1 vssd1 vccd1 vccd1 _26235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23447_ _23624_/A vssd1 vssd1 vccd1 vccd1 _23447_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20659_ _20659_/A vssd1 vssd1 vccd1 vccd1 _20659_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _13200_/A vssd1 vssd1 vccd1 vccd1 _27041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14180_ _26736_/Q _14173_/X _14167_/X _14179_/Y vssd1 vssd1 vccd1 vccd1 _26736_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26166_ _19891_/X _26166_/D vssd1 vssd1 vccd1 vccd1 _26166_/Q sky130_fd_sc_hd__dfxtp_1
X_23378_ _27765_/Q vssd1 vssd1 vccd1 vccd1 _24877_/A sky130_fd_sc_hd__buf_2
XFILLER_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13131_ _27289_/Q _13142_/B vssd1 vssd1 vccd1 vccd1 _13131_/X sky130_fd_sc_hd__and2_2
X_25117_ _25143_/A vssd1 vssd1 vccd1 vccd1 _25139_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22329_ _22315_/X _22316_/X _22317_/X _22318_/X _22319_/X _22320_/X vssd1 vssd1 vccd1
+ vccd1 _22330_/A sky130_fd_sc_hd__mux4_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26097_ _19653_/X _26097_/D vssd1 vssd1 vccd1 vccd1 _26097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25048_ _25046_/X _25047_/X _25074_/S vssd1 vssd1 vccd1 vccd1 _25048_/X sky130_fd_sc_hd__mux2_1
X_13062_ _13062_/A vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_180_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17870_ _18182_/A vssd1 vssd1 vccd1 vccd1 _17870_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16821_ _16815_/X _16820_/X _16806_/X vssd1 vssd1 vccd1 vccd1 _16821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26999_ _22800_/X _26999_/D vssd1 vssd1 vccd1 vccd1 _26999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19540_ _19534_/X _19536_/X _19539_/X _18837_/X _19312_/S vssd1 vssd1 vccd1 vccd1
+ _19549_/B sky130_fd_sc_hd__a221o_1
XFILLER_24_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16752_ _16752_/A _16752_/B vssd1 vssd1 vccd1 vccd1 _16753_/A sky130_fd_sc_hd__xor2_1
X_13964_ _13964_/A vssd1 vssd1 vccd1 vccd1 _14038_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15703_ _15703_/A _15703_/B vssd1 vssd1 vccd1 vccd1 _15703_/Y sky130_fd_sc_hd__nor2_1
X_19471_ _19471_/A _19471_/B _19471_/C vssd1 vssd1 vccd1 vccd1 _19472_/A sky130_fd_sc_hd__and3_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16683_ _16678_/Y _16679_/X _16681_/X _16682_/X vssd1 vssd1 vccd1 vccd1 _24226_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_13895_ _13895_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18422_ _18415_/X _18417_/X _18421_/X _18285_/X _18372_/X vssd1 vssd1 vccd1 vccd1
+ _18423_/C sky130_fd_sc_hd__a221o_1
X_15634_ _13078_/X _26165_/Q _15634_/S vssd1 vssd1 vccd1 vccd1 _15635_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _19313_/A _18353_/B vssd1 vssd1 vccd1 vccd1 _18354_/A sky130_fd_sc_hd__and2_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _26196_/Q _14727_/A _15573_/S vssd1 vssd1 vccd1 vccd1 _15566_/A sky130_fd_sc_hd__mux2_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17304_ _25835_/Q _26034_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17304_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14516_ _15769_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14516_/Y sky130_fd_sc_hd__nor2_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18284_ _18282_/X _18283_/X _18331_/S vssd1 vssd1 vccd1 vccd1 _18284_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15496_ _15496_/A vssd1 vssd1 vccd1 vccd1 _26227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17235_ _17233_/X _17234_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17235_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14447_ _26642_/Q _14441_/X _14437_/X _14446_/Y vssd1 vssd1 vccd1 vccd1 _26642_/D
+ sky130_fd_sc_hd__a31o_1
X_17166_ _27839_/Q _27143_/Q _25888_/Q _25856_/Q _17142_/X _17130_/X vssd1 vssd1 vccd1
+ vccd1 _17166_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14378_ _14548_/A vssd1 vssd1 vccd1 vccd1 _14441_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _16233_/C vssd1 vssd1 vccd1 vccd1 _16274_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_7_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13329_ _26999_/Q _13328_/X _13335_/S vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17097_ _25818_/Q _26017_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17097_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16048_ _27478_/Q _27374_/Q vssd1 vssd1 vccd1 vccd1 _16048_/X sky130_fd_sc_hd__and2_1
XFILLER_142_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19807_ _19807_/A vssd1 vssd1 vccd1 vccd1 _19807_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17999_ _18462_/A vssd1 vssd1 vccd1 vccd1 _17999_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19738_ _19726_/X _19727_/X _19728_/X _19729_/X _19731_/X _19733_/X vssd1 vssd1 vccd1
+ vccd1 _19739_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19669_ _19669_/A vssd1 vssd1 vccd1 vccd1 _19669_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21700_ _21700_/A vssd1 vssd1 vccd1 vccd1 _21700_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22680_ _22680_/A vssd1 vssd1 vccd1 vccd1 _22680_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21631_ _21647_/A vssd1 vssd1 vccd1 vccd1 _21631_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24350_ _27558_/Q _24350_/B vssd1 vssd1 vccd1 vccd1 _24351_/A sky130_fd_sc_hd__and2_1
X_21562_ _21562_/A vssd1 vssd1 vccd1 vccd1 _21562_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23301_ input61/X vssd1 vssd1 vccd1 vccd1 _23301_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20513_ _20513_/A vssd1 vssd1 vccd1 vccd1 _20513_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21493_ _21579_/A vssd1 vssd1 vccd1 vccd1 _21561_/A sky130_fd_sc_hd__clkbuf_2
X_24281_ _16233_/X _16234_/X _16235_/X _24279_/X vssd1 vssd1 vccd1 vccd1 _27417_/D
+ sky130_fd_sc_hd__o31a_2
XFILLER_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26020_ _26020_/CLK _26020_/D vssd1 vssd1 vccd1 vccd1 _26020_/Q sky130_fd_sc_hd__dfxtp_1
X_23232_ _23232_/A vssd1 vssd1 vccd1 vccd1 _27151_/D sky130_fd_sc_hd__clkbuf_1
X_20444_ _20702_/A vssd1 vssd1 vccd1 vccd1 _20512_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23163_ _27121_/Q _17750_/X _23165_/S vssd1 vssd1 vccd1 vccd1 _23164_/A sky130_fd_sc_hd__mux2_1
X_20375_ _20375_/A vssd1 vssd1 vccd1 vccd1 _20375_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22114_ _22162_/A vssd1 vssd1 vccd1 vccd1 _22114_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23094_ _23094_/A vssd1 vssd1 vccd1 vccd1 _23103_/S sky130_fd_sc_hd__buf_2
XFILLER_133_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27971_ _27971_/A _15940_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
X_22045_ _22035_/X _22036_/X _22037_/X _22038_/X _22039_/X _22040_/X vssd1 vssd1 vccd1
+ vccd1 _22046_/A sky130_fd_sc_hd__mux4_1
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26922_ _22532_/X _26922_/D vssd1 vssd1 vccd1 vccd1 _26922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_625 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26853_ _22296_/X _26853_/D vssd1 vssd1 vccd1 vccd1 _26853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25804_ _25804_/A vssd1 vssd1 vccd1 vccd1 _27856_/D sky130_fd_sc_hd__clkbuf_1
X_26784_ _22050_/X _26784_/D vssd1 vssd1 vccd1 vccd1 _26784_/Q sky130_fd_sc_hd__dfxtp_1
X_23996_ _23992_/X _23994_/X _24031_/S vssd1 vssd1 vccd1 vccd1 _23996_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25735_ _27379_/Q _25735_/B _25735_/C vssd1 vssd1 vccd1 vccd1 _25792_/A sky130_fd_sc_hd__or3_4
X_22947_ _22939_/X _22940_/X _22941_/X _22942_/X _22943_/X _22944_/X vssd1 vssd1 vccd1
+ vccd1 _22948_/A sky130_fd_sc_hd__mux4_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13680_ _13859_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13680_/Y sky130_fd_sc_hd__nor2_1
X_25666_ _25666_/A vssd1 vssd1 vccd1 vccd1 _25666_/X sky130_fd_sc_hd__clkbuf_1
X_22878_ _22878_/A vssd1 vssd1 vccd1 vccd1 _22878_/X sky130_fd_sc_hd__clkbuf_1
X_27405_ _27406_/CLK _27405_/D vssd1 vssd1 vccd1 vccd1 _27405_/Q sky130_fd_sc_hd__dfxtp_1
X_24617_ _24617_/A vssd1 vssd1 vccd1 vccd1 _27567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21829_ _22087_/A vssd1 vssd1 vccd1 vccd1 _21899_/A sky130_fd_sc_hd__buf_2
X_25597_ _24806_/A _25564_/X _25595_/X _25596_/Y _25592_/X vssd1 vssd1 vccd1 vccd1
+ _27780_/D sky130_fd_sc_hd__a221oi_1
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15350_ _15350_/A vssd1 vssd1 vccd1 vccd1 _26292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27336_ _27338_/CLK _27336_/D vssd1 vssd1 vccd1 vccd1 _27336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24548_ _24534_/X _24394_/A _24551_/S vssd1 vssd1 vccd1 vccd1 _24549_/B sky130_fd_sc_hd__mux2_1
XFILLER_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ _26692_/Q _14296_/X _14297_/X _14300_/Y vssd1 vssd1 vccd1 vccd1 _26692_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15281_ _15281_/A vssd1 vssd1 vccd1 vccd1 _26322_/D sky130_fd_sc_hd__clkbuf_1
X_27267_ _27335_/CLK _27267_/D vssd1 vssd1 vccd1 vccd1 _27267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24479_ _24479_/A vssd1 vssd1 vccd1 vccd1 _27515_/D sky130_fd_sc_hd__clkbuf_1
X_17020_ _16992_/X _17020_/B vssd1 vssd1 vccd1 vccd1 _17020_/X sky130_fd_sc_hd__and2b_1
X_14232_ _14410_/A _14234_/B vssd1 vssd1 vccd1 vccd1 _14232_/Y sky130_fd_sc_hd__nor2_1
X_26218_ _20073_/X _26218_/D vssd1 vssd1 vccd1 vccd1 _26218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27198_ _27209_/CLK _27198_/D vssd1 vssd1 vccd1 vccd1 _27198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ _26742_/Q _14157_/X _14151_/X _14162_/Y vssd1 vssd1 vccd1 vccd1 _26742_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_124_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26149_ _19829_/X _26149_/D vssd1 vssd1 vccd1 vccd1 _26149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ _27292_/Q _13142_/B vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__and2_2
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14094_ _14359_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14094_/Y sky130_fd_sc_hd__nor2_1
X_18971_ _18775_/X _18970_/X _18941_/X vssd1 vssd1 vccd1 vccd1 _18971_/X sky130_fd_sc_hd__o21a_1
XFILLER_125_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _18403_/A vssd1 vssd1 vccd1 vccd1 _17922_/X sky130_fd_sc_hd__clkbuf_4
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13045_ _27267_/Q vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17853_ _18443_/A vssd1 vssd1 vccd1 vccd1 _18285_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16804_ _16804_/A _16804_/B vssd1 vssd1 vccd1 vccd1 _16804_/Y sky130_fd_sc_hd__nor2_1
X_14996_ _15023_/A vssd1 vssd1 vccd1 vccd1 _15008_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17784_ _18455_/A vssd1 vssd1 vccd1 vccd1 _18481_/A sky130_fd_sc_hd__buf_4
XFILLER_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19523_ _26167_/Q _26103_/Q _27031_/Q _26999_/Q _19460_/X _19482_/X vssd1 vssd1 vccd1
+ vccd1 _19524_/B sky130_fd_sc_hd__mux4_1
X_13947_ _14331_/A _13954_/B vssd1 vssd1 vccd1 vccd1 _13947_/Y sky130_fd_sc_hd__nor2_1
X_16735_ _16084_/A _16733_/X _16734_/X vssd1 vssd1 vccd1 vccd1 _16735_/X sky130_fd_sc_hd__o21ba_1
X_19454_ _26708_/Q _26676_/Q _26644_/Q _26612_/Q _18816_/X _19385_/X vssd1 vssd1 vccd1
+ vccd1 _19454_/X sky130_fd_sc_hd__mux4_1
X_16666_ _16816_/A _16666_/B vssd1 vssd1 vccd1 vccd1 _16666_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_24 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13878_ _13878_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18405_ _18405_/A vssd1 vssd1 vccd1 vccd1 _18532_/S sky130_fd_sc_hd__clkbuf_2
X_15617_ _26172_/Q _14804_/A _15617_/S vssd1 vssd1 vccd1 vccd1 _15618_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19385_ _19385_/A vssd1 vssd1 vccd1 vccd1 _19385_/X sky130_fd_sc_hd__clkbuf_2
X_16597_ _16599_/A _16599_/B vssd1 vssd1 vccd1 vccd1 _16878_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18336_ _18336_/A _18379_/A vssd1 vssd1 vccd1 vccd1 _18336_/X sky130_fd_sc_hd__or2b_1
X_15548_ _15548_/A vssd1 vssd1 vccd1 vccd1 _26203_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18267_ _18425_/A vssd1 vssd1 vccd1 vccd1 _18267_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15479_ _15783_/B _15551_/B vssd1 vssd1 vccd1 vccd1 _15536_/A sky130_fd_sc_hd__or2_2
XFILLER_129_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17218_ _17216_/X _17218_/B vssd1 vssd1 vccd1 vccd1 _17218_/X sky130_fd_sc_hd__and2b_1
XFILLER_147_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18198_ _18379_/A vssd1 vssd1 vccd1 vccd1 _18198_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17149_ _17116_/X _17143_/X _17146_/X _17148_/X vssd1 vssd1 vccd1 vccd1 _17149_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20160_ _20146_/X _20147_/X _20148_/X _20149_/X _20150_/X _20151_/X vssd1 vssd1 vccd1
+ vccd1 _20161_/A sky130_fd_sc_hd__mux4_1
XFILLER_144_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20091_ _20091_/A vssd1 vssd1 vccd1 vccd1 _20091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23850_ _23991_/A vssd1 vssd1 vccd1 vccd1 _23850_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22801_ _22887_/A vssd1 vssd1 vccd1 vccd1 _22869_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23781_ _27068_/Q _27100_/Q _23796_/S vssd1 vssd1 vccd1 vccd1 _23781_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20993_ _21041_/A vssd1 vssd1 vccd1 vccd1 _20993_/X sky130_fd_sc_hd__clkbuf_1
X_25520_ _24769_/A _25504_/X _25516_/Y _25519_/X _25497_/X vssd1 vssd1 vccd1 vccd1
+ _27767_/D sky130_fd_sc_hd__a221oi_1
XFILLER_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22732_ _22732_/A vssd1 vssd1 vccd1 vccd1 _22732_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25451_ _24267_/A _25440_/X _25442_/X _24832_/B _24384_/A vssd1 vssd1 vccd1 vccd1
+ _25451_/X sky130_fd_sc_hd__o311a_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22663_ _22649_/X _22650_/X _22651_/X _22652_/X _22653_/X _22654_/X vssd1 vssd1 vccd1
+ vccd1 _22664_/A sky130_fd_sc_hd__mux4_1
XFILLER_201_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24402_ _24538_/A vssd1 vssd1 vccd1 vccd1 _24411_/B sky130_fd_sc_hd__clkbuf_1
X_21614_ _21614_/A vssd1 vssd1 vccd1 vccd1 _21614_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25382_ _25428_/S vssd1 vssd1 vccd1 vccd1 _25391_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_200_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22594_ _22610_/A vssd1 vssd1 vccd1 vccd1 _22594_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27121_ _27121_/CLK _27121_/D vssd1 vssd1 vccd1 vccd1 _27121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24333_ _27550_/Q _24339_/B vssd1 vssd1 vccd1 vccd1 _24334_/A sky130_fd_sc_hd__and2_1
X_21545_ _21561_/A vssd1 vssd1 vccd1 vccd1 _21545_/X sky130_fd_sc_hd__clkbuf_1
X_27052_ _22988_/X _27052_/D vssd1 vssd1 vccd1 vccd1 _27052_/Q sky130_fd_sc_hd__dfxtp_1
X_24264_ _24264_/A _24264_/B vssd1 vssd1 vccd1 vccd1 _27406_/D sky130_fd_sc_hd__nor2_1
X_21476_ _21476_/A vssd1 vssd1 vccd1 vccd1 _21476_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26003_ _27092_/CLK _26003_/D vssd1 vssd1 vccd1 vccd1 _26003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23215_ _17469_/X _27144_/Q _23215_/S vssd1 vssd1 vccd1 vccd1 _23216_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20427_ _20427_/A vssd1 vssd1 vccd1 vccd1 _20427_/X sky130_fd_sc_hd__clkbuf_1
X_24195_ _27473_/Q _24195_/B vssd1 vssd1 vccd1 vccd1 _24196_/A sky130_fd_sc_hd__and2_1
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23146_ _27113_/Q _17724_/X _23154_/S vssd1 vssd1 vccd1 vccd1 _23147_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20358_ _25657_/A vssd1 vssd1 vccd1 vccd1 _20706_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23077_ _27083_/Q _17731_/X _23081_/S vssd1 vssd1 vccd1 vccd1 _23078_/A sky130_fd_sc_hd__mux2_1
X_27954_ _27954_/A _15921_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
XFILLER_122_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20289_ _20337_/A vssd1 vssd1 vccd1 vccd1 _20289_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22028_ _22028_/A vssd1 vssd1 vccd1 vccd1 _22028_/X sky130_fd_sc_hd__clkbuf_1
X_26905_ _22478_/X _26905_/D vssd1 vssd1 vccd1 vccd1 _26905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14850_ _14850_/A vssd1 vssd1 vccd1 vccd1 _26506_/D sky130_fd_sc_hd__clkbuf_1
X_26836_ _22238_/X _26836_/D vssd1 vssd1 vccd1 vccd1 _26836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13801_ _13827_/A vssd1 vssd1 vccd1 vccd1 _13812_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_26767_ _21992_/X _26767_/D vssd1 vssd1 vccd1 vccd1 _26767_/Q sky130_fd_sc_hd__dfxtp_1
X_14781_ _14781_/A vssd1 vssd1 vccd1 vccd1 _26532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23979_ _27089_/Q _27121_/Q _23986_/S vssd1 vssd1 vccd1 vccd1 _23979_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16520_ _16824_/B _16550_/B vssd1 vssd1 vccd1 vccd1 _16662_/A sky130_fd_sc_hd__xnor2_1
X_13732_ _13745_/A vssd1 vssd1 vccd1 vccd1 _13732_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25718_ _25718_/A vssd1 vssd1 vccd1 vccd1 _25718_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26698_ _21754_/X _26698_/D vssd1 vssd1 vccd1 vccd1 _26698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16451_ _16451_/A _16563_/B vssd1 vssd1 vccd1 vccd1 _16451_/Y sky130_fd_sc_hd__nor2_1
X_13663_ _13934_/A _13670_/B vssd1 vssd1 vccd1 vccd1 _13663_/Y sky130_fd_sc_hd__nor2_1
X_25649_ _25635_/X _25636_/X _25637_/X _25638_/X _25640_/X _25642_/X vssd1 vssd1 vccd1
+ vccd1 _25650_/A sky130_fd_sc_hd__mux4_1
XFILLER_188_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15402_ _15402_/A vssd1 vssd1 vccd1 vccd1 _26268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19343_/A vssd1 vssd1 vccd1 vccd1 _19170_/X sky130_fd_sc_hd__buf_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _16751_/B _16398_/B vssd1 vssd1 vccd1 vccd1 _16383_/B sky130_fd_sc_hd__nand2_1
X_13594_ _26935_/Q _13580_/X _13587_/X _13593_/Y vssd1 vssd1 vccd1 vccd1 _26935_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _18118_/X _18119_/X _18216_/S vssd1 vssd1 vccd1 vccd1 _18121_/X sky130_fd_sc_hd__mux2_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15333_ _15333_/A vssd1 vssd1 vccd1 vccd1 _26298_/D sky130_fd_sc_hd__clkbuf_1
X_27319_ _27328_/CLK _27319_/D vssd1 vssd1 vccd1 vccd1 _27319_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18052_ _18146_/A _18052_/B _18052_/C vssd1 vssd1 vccd1 vccd1 _18053_/A sky130_fd_sc_hd__and3_1
X_15264_ _15332_/S vssd1 vssd1 vccd1 vccd1 _15273_/S sky130_fd_sc_hd__buf_2
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17003_ _16985_/X _16990_/X _16996_/X _17002_/X vssd1 vssd1 vccd1 vccd1 _17003_/X
+ sky130_fd_sc_hd__o22a_1
X_14215_ _14215_/A vssd1 vssd1 vccd1 vccd1 _14226_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_5 _21442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15195_ _14715_/X _26360_/Q _15201_/S vssd1 vssd1 vccd1 vccd1 _15196_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _26747_/Q _14142_/X _14070_/B _14145_/Y vssd1 vssd1 vccd1 vccd1 _26747_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_113_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14077_ _14342_/A _14085_/B vssd1 vssd1 vccd1 vccd1 _14077_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18954_ _19485_/A vssd1 vssd1 vccd1 vccd1 _18954_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17905_ _26396_/Q _26364_/Q _26332_/Q _26300_/Q _17903_/X _17904_/X vssd1 vssd1 vccd1
+ vccd1 _17905_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13028_ _13102_/A vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__clkbuf_4
X_18885_ _26268_/Q _26236_/Q _26204_/Q _26172_/Q _18859_/X _18818_/X vssd1 vssd1 vccd1
+ vccd1 _18885_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17836_ _26266_/Q _26234_/Q _26202_/Q _26170_/Q _17832_/X _17835_/X vssd1 vssd1 vccd1
+ vccd1 _17836_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17767_ _25940_/Q _17766_/X _17770_/S vssd1 vssd1 vccd1 vccd1 _17768_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14979_ _15716_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14979_/Y sky130_fd_sc_hd__nor2_1
X_19506_ _19524_/A _19506_/B vssd1 vssd1 vccd1 vccd1 _19506_/X sky130_fd_sc_hd__or2_1
X_16718_ _16719_/A _16719_/B _16719_/C vssd1 vssd1 vccd1 vccd1 _16890_/C sky130_fd_sc_hd__a21o_1
X_17698_ _17698_/A vssd1 vssd1 vccd1 vccd1 _25918_/D sky130_fd_sc_hd__clkbuf_1
X_19437_ _19430_/X _19433_/X _19436_/X _19324_/X _19393_/X vssd1 vssd1 vccd1 vccd1
+ _19450_/B sky130_fd_sc_hd__a221o_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16649_ _16623_/A _16648_/B _16648_/C vssd1 vssd1 vccd1 vccd1 _16650_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19368_ _26704_/Q _26672_/Q _26640_/Q _26608_/Q _18767_/X _18909_/X vssd1 vssd1 vccd1
+ vccd1 _19369_/B sky130_fd_sc_hd__mux4_2
XFILLER_124_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18319_ _18198_/X _18315_/X _18318_/X _18203_/X vssd1 vssd1 vccd1 vccd1 _18319_/X
+ sky130_fd_sc_hd__o211a_1
X_19299_ _19299_/A _19299_/B vssd1 vssd1 vccd1 vccd1 _19299_/X sky130_fd_sc_hd__or2_1
XFILLER_191_802 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21330_ _21378_/A vssd1 vssd1 vccd1 vccd1 _21330_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21261_ _21253_/X _21254_/X _21255_/X _21256_/X _21257_/X _21258_/X vssd1 vssd1 vccd1
+ vccd1 _21262_/A sky130_fd_sc_hd__mux4_1
X_23000_ _23000_/A vssd1 vssd1 vccd1 vccd1 _23000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20212_ _20200_/X _20201_/X _20202_/X _20203_/X _20204_/X _20205_/X vssd1 vssd1 vccd1
+ vccd1 _20213_/A sky130_fd_sc_hd__mux4_1
X_21192_ _21192_/A vssd1 vssd1 vccd1 vccd1 _21192_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20143_ _20143_/A vssd1 vssd1 vccd1 vccd1 _20143_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20074_ _20060_/X _20061_/X _20062_/X _20063_/X _20064_/X _20065_/X vssd1 vssd1 vccd1
+ vccd1 _20075_/A sky130_fd_sc_hd__mux4_1
X_24951_ _24954_/B _24954_/C vssd1 vssd1 vccd1 vccd1 _24952_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23902_ _23898_/X _23900_/X _23938_/S vssd1 vssd1 vccd1 vccd1 _23902_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27670_ _27754_/CLK _27670_/D vssd1 vssd1 vccd1 vccd1 _27670_/Q sky130_fd_sc_hd__dfxtp_1
X_24882_ _24887_/B _24882_/B vssd1 vssd1 vccd1 vccd1 _24883_/B sky130_fd_sc_hd__or2_1
XFILLER_44_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater350 _27754_/CLK vssd1 vssd1 vccd1 vccd1 _27645_/CLK sky130_fd_sc_hd__clkbuf_1
X_26621_ _21486_/X _26621_/D vssd1 vssd1 vccd1 vccd1 _26621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater361 _25909_/CLK vssd1 vssd1 vccd1 vccd1 _27572_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater372 _27342_/CLK vssd1 vssd1 vccd1 vccd1 _27682_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23833_ _23800_/X _23831_/X _23832_/X _23816_/X vssd1 vssd1 vccd1 vccd1 _27278_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater383 _27207_/CLK vssd1 vssd1 vccd1 vccd1 _27450_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater394 _27825_/CLK vssd1 vssd1 vccd1 vccd1 _27341_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26552_ _21248_/X _26552_/D vssd1 vssd1 vccd1 vccd1 _26552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23764_ _24003_/A vssd1 vssd1 vccd1 vccd1 _23862_/A sky130_fd_sc_hd__buf_2
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _21041_/A vssd1 vssd1 vccd1 vccd1 _20976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25503_ _24763_/A _25474_/X _25499_/Y _25502_/X _25497_/X vssd1 vssd1 vccd1 vccd1
+ _27764_/D sky130_fd_sc_hd__a221oi_1
XFILLER_14_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22715_ _22887_/A vssd1 vssd1 vccd1 vccd1 _22783_/A sky130_fd_sc_hd__buf_2
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26483_ _21004_/X _26483_/D vssd1 vssd1 vccd1 vccd1 _26483_/Q sky130_fd_sc_hd__dfxtp_1
X_23695_ _23695_/A vssd1 vssd1 vccd1 vccd1 _27252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25434_ _25434_/A vssd1 vssd1 vccd1 vccd1 _25569_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_198_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22646_ _22646_/A vssd1 vssd1 vccd1 vccd1 _22646_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25365_ _27723_/Q input63/X _25369_/S vssd1 vssd1 vccd1 vccd1 _25366_/A sky130_fd_sc_hd__mux2_1
X_22577_ _22609_/A vssd1 vssd1 vccd1 vccd1 _22577_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27104_ _27105_/CLK _27104_/D vssd1 vssd1 vccd1 vccd1 _27104_/Q sky130_fd_sc_hd__dfxtp_1
X_24316_ _24316_/A vssd1 vssd1 vccd1 vccd1 _27442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21528_ _21528_/A vssd1 vssd1 vccd1 vccd1 _21528_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25296_ _25306_/A _25296_/B vssd1 vssd1 vccd1 vccd1 _25296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27035_ _22930_/X _27035_/D vssd1 vssd1 vccd1 vccd1 _27035_/Q sky130_fd_sc_hd__dfxtp_1
X_24247_ _24247_/A _24250_/B vssd1 vssd1 vccd1 vccd1 _24248_/A sky130_fd_sc_hd__and2_1
X_21459_ _21475_/A vssd1 vssd1 vccd1 vccd1 _21459_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14000_ _26795_/Q _13987_/X _13983_/X _13999_/Y vssd1 vssd1 vccd1 vccd1 _26795_/D
+ sky130_fd_sc_hd__a31o_1
X_24178_ _27465_/Q _24184_/B vssd1 vssd1 vccd1 vccd1 _24179_/A sky130_fd_sc_hd__and2_1
XFILLER_123_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23129_ _23129_/A vssd1 vssd1 vccd1 vccd1 _27105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15951_ _15955_/A vssd1 vssd1 vccd1 vccd1 _15951_/Y sky130_fd_sc_hd__inv_2
X_27937_ _27937_/A _15946_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14902_ _14902_/A vssd1 vssd1 vccd1 vccd1 _26483_/D sky130_fd_sc_hd__clkbuf_1
X_18670_ _26000_/Q _17747_/X _18674_/S vssd1 vssd1 vccd1 vccd1 _18671_/A sky130_fd_sc_hd__mux2_1
X_15882_ _15894_/A vssd1 vssd1 vccd1 vccd1 _15887_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17621_ _17450_/X _25883_/Q _17623_/S vssd1 vssd1 vccd1 vccd1 _17622_/A sky130_fd_sc_hd__mux2_1
X_26819_ _22172_/X _26819_/D vssd1 vssd1 vccd1 vccd1 _26819_/Q sky130_fd_sc_hd__dfxtp_1
X_14833_ _26513_/Q _13347_/X _14835_/S vssd1 vssd1 vccd1 vccd1 _14834_/A sky130_fd_sc_hd__mux2_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27799_ _25648_/X _27799_/D vssd1 vssd1 vccd1 vccd1 _27799_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _17552_/A vssd1 vssd1 vccd1 vccd1 _25852_/D sky130_fd_sc_hd__clkbuf_1
X_14764_ _14763_/X _26537_/Q _14773_/S vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__mux2_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13715_ _26892_/Q _13710_/X _13705_/X _13714_/Y vssd1 vssd1 vccd1 vccd1 _26892_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16503_ _14750_/A _16501_/X _16311_/X _25963_/Q _16502_/Y vssd1 vssd1 vccd1 vccd1
+ _16632_/B sky130_fd_sc_hd__a221o_1
XFILLER_60_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17483_ _17482_/X _25829_/Q _17486_/S vssd1 vssd1 vccd1 vccd1 _17484_/A sky130_fd_sc_hd__mux2_1
X_14695_ _26560_/Q _14685_/X _14693_/X _14694_/Y vssd1 vssd1 vccd1 vccd1 _26560_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19222_ _19222_/A _19222_/B _19222_/C vssd1 vssd1 vccd1 vccd1 _19223_/A sky130_fd_sc_hd__and3_1
X_13646_ _26916_/Q _13639_/X _13642_/X _13645_/Y vssd1 vssd1 vccd1 vccd1 _26916_/D
+ sky130_fd_sc_hd__a31o_1
X_16434_ _14769_/A _16384_/X _16412_/A _25957_/Q vssd1 vssd1 vccd1 vccd1 _16434_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _27381_/Q _16402_/A vssd1 vssd1 vccd1 vccd1 _16365_/Y sky130_fd_sc_hd__nand2_1
X_19153_ _19222_/A _19153_/B _19153_/C vssd1 vssd1 vccd1 vccd1 _19154_/A sky130_fd_sc_hd__and3_1
X_13577_ _13938_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13577_/Y sky130_fd_sc_hd__nor2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18104_ _18100_/X _18102_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18104_/X sky130_fd_sc_hd__mux2_1
X_15316_ _15316_/A vssd1 vssd1 vccd1 vccd1 _26306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16296_ _16298_/B _16296_/B _26067_/Q vssd1 vssd1 vccd1 vccd1 _16296_/X sky130_fd_sc_hd__or3b_2
XFILLER_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19084_ _19084_/A vssd1 vssd1 vccd1 vccd1 _26051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18035_ _26817_/Q _26785_/Q _26753_/Q _26721_/Q _18034_/X _17890_/X vssd1 vssd1 vccd1
+ vccd1 _18035_/X sky130_fd_sc_hd__mux4_1
X_15247_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15256_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_172_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15178_ _26367_/Q _13405_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14129_ _26754_/Q _14117_/X _14120_/X _14128_/Y vssd1 vssd1 vccd1 vccd1 _26754_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19986_ _19972_/X _19973_/X _19974_/X _19975_/X _19976_/X _19977_/X vssd1 vssd1 vccd1
+ vccd1 _19987_/A sky130_fd_sc_hd__mux4_1
XFILLER_154_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18937_ _26814_/Q _26782_/Q _26750_/Q _26718_/Q _18870_/X _18770_/X vssd1 vssd1 vccd1
+ vccd1 _18938_/B sky130_fd_sc_hd__mux4_1
XFILLER_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18868_ _18989_/A _18868_/B _18868_/C vssd1 vssd1 vccd1 vccd1 _18869_/A sky130_fd_sc_hd__and3_1
X_17819_ _18412_/A vssd1 vssd1 vccd1 vccd1 _24396_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18799_ _18791_/X _18796_/X _19560_/A vssd1 vssd1 vccd1 vccd1 _18799_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20830_ _20816_/X _20817_/X _20818_/X _20819_/X _20820_/X _20821_/X vssd1 vssd1 vccd1
+ vccd1 _20831_/A sky130_fd_sc_hd__mux4_1
XFILLER_82_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20761_ _20761_/A vssd1 vssd1 vccd1 vccd1 _20761_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22500_ _22500_/A vssd1 vssd1 vccd1 vccd1 _22500_/X sky130_fd_sc_hd__clkbuf_1
X_23480_ _27185_/Q _23483_/B vssd1 vssd1 vccd1 vccd1 _23480_/X sky130_fd_sc_hd__or2_1
XFILLER_196_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20692_ _20684_/X _20685_/X _20686_/X _20687_/X _20689_/X _20691_/X vssd1 vssd1 vccd1
+ vccd1 _20693_/A sky130_fd_sc_hd__mux4_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22431_ _22417_/X _22418_/X _22419_/X _22420_/X _22421_/X _22422_/X vssd1 vssd1 vccd1
+ vccd1 _22432_/A sky130_fd_sc_hd__mux4_1
XFILLER_202_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25150_ _25150_/A _25150_/B vssd1 vssd1 vccd1 vccd1 _25151_/B sky130_fd_sc_hd__xnor2_1
XFILLER_175_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22362_ _22362_/A vssd1 vssd1 vccd1 vccd1 _22362_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24101_ _24101_/A vssd1 vssd1 vccd1 vccd1 _27325_/D sky130_fd_sc_hd__clkbuf_1
X_21313_ _21301_/X _21302_/X _21303_/X _21304_/X _21307_/X _21310_/X vssd1 vssd1 vccd1
+ vccd1 _21314_/A sky130_fd_sc_hd__mux4_1
X_25081_ _27078_/Q _27110_/Q _25088_/S vssd1 vssd1 vccd1 vccd1 _25081_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22293_ _22280_/X _22282_/X _22284_/X _22286_/X _22287_/X _22288_/X vssd1 vssd1 vccd1
+ vccd1 _22294_/A sky130_fd_sc_hd__mux4_1
X_24032_ _27095_/Q _27127_/Q _24032_/S vssd1 vssd1 vccd1 vccd1 _24032_/X sky130_fd_sc_hd__mux2_1
X_21244_ _21244_/A vssd1 vssd1 vccd1 vccd1 _21244_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21175_ _21163_/X _21164_/X _21165_/X _21166_/X _21167_/X _21168_/X vssd1 vssd1 vccd1
+ vccd1 _21176_/A sky130_fd_sc_hd__mux4_1
XFILLER_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20126_ _20114_/X _20115_/X _20116_/X _20117_/X _20118_/X _20119_/X vssd1 vssd1 vccd1
+ vccd1 _20127_/A sky130_fd_sc_hd__mux4_1
X_25983_ _26016_/CLK _25983_/D vssd1 vssd1 vccd1 vccd1 _25983_/Q sky130_fd_sc_hd__dfxtp_1
X_20057_ _20057_/A vssd1 vssd1 vccd1 vccd1 _20057_/X sky130_fd_sc_hd__clkbuf_1
X_27722_ _27750_/CLK _27722_/D vssd1 vssd1 vccd1 vccd1 _27722_/Q sky130_fd_sc_hd__dfxtp_1
X_24934_ _27663_/Q _24909_/X _24933_/Y _24914_/X vssd1 vssd1 vccd1 vccd1 _27663_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27653_ _27654_/CLK _27653_/D vssd1 vssd1 vccd1 vccd1 _27653_/Q sky130_fd_sc_hd__dfxtp_1
X_24865_ _27649_/Q _24861_/X _24863_/Y _24864_/X vssd1 vssd1 vccd1 vccd1 _27649_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater180 _27674_/CLK vssd1 vssd1 vccd1 vccd1 _27096_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater191 _25980_/CLK vssd1 vssd1 vccd1 vccd1 _26016_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_203 _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26604_ _21426_/X _26604_/D vssd1 vssd1 vccd1 vccd1 _26604_/Q sky130_fd_sc_hd__dfxtp_1
X_23816_ _23864_/A vssd1 vssd1 vccd1 vccd1 _23816_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _14518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27584_ _27584_/CLK _27584_/D vssd1 vssd1 vccd1 vccd1 _27584_/Q sky130_fd_sc_hd__dfxtp_1
X_24796_ _24796_/A _24800_/B vssd1 vssd1 vccd1 vccd1 _24796_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_225 _14810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_236 _17321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _27772_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26535_ _21186_/X _26535_/D vssd1 vssd1 vccd1 vccd1 _26535_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_258 _26816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23747_ _23946_/A vssd1 vssd1 vccd1 vccd1 _23747_/X sky130_fd_sc_hd__buf_2
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20959_ _21217_/A vssd1 vssd1 vccd1 vccd1 _21028_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_187_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13500_ _26956_/Q _13487_/X _13482_/X _13499_/Y vssd1 vssd1 vccd1 vccd1 _26956_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14480_ _15743_/A _14483_/B vssd1 vssd1 vccd1 vccd1 _14480_/Y sky130_fd_sc_hd__nor2_1
X_26466_ _20946_/X _26466_/D vssd1 vssd1 vccd1 vccd1 _26466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23678_ _23678_/A vssd1 vssd1 vccd1 vccd1 _27244_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13431_ _16033_/A vssd1 vssd1 vccd1 vccd1 _13857_/A sky130_fd_sc_hd__clkbuf_2
X_25417_ _25417_/A vssd1 vssd1 vccd1 vccd1 _27746_/D sky130_fd_sc_hd__clkbuf_1
X_22629_ _22887_/A vssd1 vssd1 vccd1 vccd1 _22697_/A sky130_fd_sc_hd__clkbuf_4
X_26397_ _20697_/X _26397_/D vssd1 vssd1 vccd1 vccd1 _26397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16150_ _16148_/Y _16119_/X _16121_/X _14448_/A _16149_/Y vssd1 vssd1 vccd1 vccd1
+ _24301_/A sky130_fd_sc_hd__o221a_2
X_25348_ _25348_/A _25348_/B vssd1 vssd1 vccd1 vccd1 _25350_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13362_ _13362_/A vssd1 vssd1 vccd1 vccd1 _26989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15101_ _14788_/X _26401_/Q _15101_/S vssd1 vssd1 vccd1 vccd1 _15102_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16081_ _25911_/Q vssd1 vssd1 vccd1 vccd1 _16646_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25279_ _25332_/A vssd1 vssd1 vccd1 vccd1 _25347_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13293_ _13304_/A vssd1 vssd1 vccd1 vccd1 _13302_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_170_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15032_ _15769_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15032_/Y sky130_fd_sc_hd__nor2_1
X_27018_ _22866_/X _27018_/D vssd1 vssd1 vccd1 vccd1 _27018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19840_ _19831_/X _19833_/X _19835_/X _19837_/X _19838_/X _19839_/X vssd1 vssd1 vccd1
+ vccd1 _19841_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19771_ _19771_/A vssd1 vssd1 vccd1 vccd1 _19771_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16983_ _16983_/A vssd1 vssd1 vccd1 vccd1 _25908_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18722_ _26023_/Q _17718_/X _18724_/S vssd1 vssd1 vccd1 vccd1 _18723_/A sky130_fd_sc_hd__mux2_1
X_15934_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15934_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _18653_/A vssd1 vssd1 vccd1 vccd1 _25992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _15868_/A vssd1 vssd1 vccd1 vccd1 _15865_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _17408_/X _25875_/Q _17612_/S vssd1 vssd1 vccd1 vccd1 _17605_/A sky130_fd_sc_hd__mux2_1
X_14816_ _26521_/Q _13319_/X _14824_/S vssd1 vssd1 vccd1 vccd1 _14817_/A sky130_fd_sc_hd__mux2_1
X_18584_ _18584_/A vssd1 vssd1 vccd1 vccd1 _24828_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15796_ _15853_/S vssd1 vssd1 vccd1 vccd1 _15805_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17535_ _17535_/A vssd1 vssd1 vccd1 vccd1 _25844_/D sky130_fd_sc_hd__clkbuf_1
X_14747_ _14747_/A vssd1 vssd1 vccd1 vccd1 _14747_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_199_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17466_ _27421_/Q vssd1 vssd1 vccd1 vccd1 _17466_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14678_ _26566_/Q _14671_/X _14666_/X _14677_/Y vssd1 vssd1 vccd1 vccd1 _26566_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19205_ _19250_/A _19205_/B vssd1 vssd1 vccd1 vccd1 _19205_/X sky130_fd_sc_hd__or2_1
X_13629_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13629_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16417_ _16733_/B _16417_/B vssd1 vssd1 vccd1 vccd1 _16708_/B sky130_fd_sc_hd__xor2_2
XFILLER_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17397_ _25657_/A vssd1 vssd1 vccd1 vccd1 _19834_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater83 _27425_/CLK vssd1 vssd1 vccd1 vccd1 _27295_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater94 _26002_/CLK vssd1 vssd1 vccd1 vccd1 _27850_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19136_ _19501_/A _19136_/B vssd1 vssd1 vccd1 vccd1 _19136_/X sky130_fd_sc_hd__or2_1
X_16348_ _16864_/A _16864_/B _16347_/Y vssd1 vssd1 vccd1 vccd1 _16867_/B sky130_fd_sc_hd__a21bo_1
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19067_ _26819_/Q _26787_/Q _26755_/Q _26723_/Q _18913_/X _24400_/A vssd1 vssd1 vccd1
+ vccd1 _19067_/X sky130_fd_sc_hd__mux4_2
X_16279_ _16108_/A _16274_/X _16276_/Y _16277_/Y _16278_/X vssd1 vssd1 vccd1 vccd1
+ _16816_/A sky130_fd_sc_hd__o41a_2
XFILLER_161_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18018_ _26144_/Q _26080_/Q _27008_/Q _26976_/Q _17870_/X _17959_/X vssd1 vssd1 vccd1
+ vccd1 _18019_/A sky130_fd_sc_hd__mux4_1
XFILLER_195_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19969_ _19969_/A vssd1 vssd1 vccd1 vccd1 _19969_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22980_ _25638_/A vssd1 vssd1 vccd1 vccd1 _22980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21931_ _22017_/A vssd1 vssd1 vccd1 vccd1 _21998_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24650_ _24663_/A vssd1 vssd1 vccd1 vccd1 _24650_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21862_ _21862_/A vssd1 vssd1 vccd1 vccd1 _21862_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23601_ _24941_/A _27220_/Q _23616_/S vssd1 vssd1 vccd1 vccd1 _23602_/B sky130_fd_sc_hd__mux2_1
X_20813_ _20813_/A vssd1 vssd1 vccd1 vccd1 _20813_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24581_ _27651_/Q _24587_/B vssd1 vssd1 vccd1 vccd1 _24582_/A sky130_fd_sc_hd__and2_1
X_21793_ _21825_/A vssd1 vssd1 vccd1 vccd1 _21793_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26320_ _20435_/X _26320_/D vssd1 vssd1 vccd1 vccd1 _26320_/Q sky130_fd_sc_hd__dfxtp_1
X_23532_ _23532_/A vssd1 vssd1 vccd1 vccd1 _27200_/D sky130_fd_sc_hd__clkbuf_1
X_20744_ _20738_/X _20739_/X _20740_/X _20741_/X _20742_/X _20743_/X vssd1 vssd1 vccd1
+ vccd1 _20745_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26251_ _20193_/X _26251_/D vssd1 vssd1 vccd1 vccd1 _26251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23463_ _27178_/Q _23470_/B vssd1 vssd1 vccd1 vccd1 _23463_/X sky130_fd_sc_hd__or2_1
XFILLER_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20675_ _20675_/A vssd1 vssd1 vccd1 vccd1 _20675_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25202_ _27531_/Q _27499_/Q vssd1 vssd1 vccd1 vccd1 _25203_/B sky130_fd_sc_hd__or2_1
X_22414_ _22414_/A vssd1 vssd1 vccd1 vccd1 _22414_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26182_ _19951_/X _26182_/D vssd1 vssd1 vccd1 vccd1 _26182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23394_ _27257_/Q vssd1 vssd1 vccd1 vccd1 _23394_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25133_ _27692_/Q _25112_/X _25131_/Y _25132_/X vssd1 vssd1 vccd1 vccd1 _27692_/D
+ sky130_fd_sc_hd__o211a_1
X_22345_ _22331_/X _22332_/X _22333_/X _22334_/X _22335_/X _22336_/X vssd1 vssd1 vccd1
+ vccd1 _22346_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25064_ _25062_/X _25063_/X _25087_/S vssd1 vssd1 vccd1 vccd1 _25064_/X sky130_fd_sc_hd__mux2_1
X_22276_ _22276_/A vssd1 vssd1 vccd1 vccd1 _22276_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24015_ _27853_/Q _27157_/Q _25902_/Q _25870_/Q _24014_/X _23991_/X vssd1 vssd1 vccd1
+ vccd1 _24015_/X sky130_fd_sc_hd__mux4_1
X_21227_ _21211_/X _21212_/X _21213_/X _21214_/X _21216_/X _21218_/X vssd1 vssd1 vccd1
+ vccd1 _21228_/A sky130_fd_sc_hd__mux4_1
XFILLER_144_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21158_ _21158_/A vssd1 vssd1 vccd1 vccd1 _21158_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20109_ _20109_/A vssd1 vssd1 vccd1 vccd1 _20109_/X sky130_fd_sc_hd__clkbuf_1
X_13980_ _14452_/A vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__buf_2
XFILLER_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25966_ _17407_/Y _25966_/D vssd1 vssd1 vccd1 vccd1 _25966_/Q sky130_fd_sc_hd__dfxtp_1
X_21089_ _21077_/X _21078_/X _21079_/X _21080_/X _21081_/X _21082_/X vssd1 vssd1 vccd1
+ vccd1 _21090_/A sky130_fd_sc_hd__mux4_1
XFILLER_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27705_ _27705_/CLK _27705_/D vssd1 vssd1 vccd1 vccd1 _27705_/Q sky130_fd_sc_hd__dfxtp_1
X_12931_ input2/X _12931_/B vssd1 vssd1 vccd1 vccd1 _12932_/A sky130_fd_sc_hd__and2b_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24917_ _27773_/Q _24918_/B vssd1 vssd1 vccd1 vccd1 _24925_/C sky130_fd_sc_hd__and2_1
X_25897_ _25897_/CLK _25897_/D vssd1 vssd1 vccd1 vccd1 _25897_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27636_ _27636_/CLK _27636_/D vssd1 vssd1 vccd1 vccd1 _27636_/Q sky130_fd_sc_hd__dfxtp_1
X_15650_ _13122_/X _26158_/Q _15656_/S vssd1 vssd1 vccd1 vccd1 _15651_/A sky130_fd_sc_hd__mux2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24848_ _24848_/A _24851_/C vssd1 vssd1 vccd1 vccd1 _24849_/B sky130_fd_sc_hd__xnor2_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _26594_/Q _14589_/X _14592_/X _14600_/Y vssd1 vssd1 vccd1 vccd1 _26594_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15581_/A vssd1 vssd1 vccd1 vccd1 _26189_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24779_ _27625_/Q _24771_/X _24778_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _27625_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27567_ _27569_/CLK _27567_/D vssd1 vssd1 vccd1 vccd1 _27567_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _27091_/Q _27123_/Q _17355_/S vssd1 vssd1 vccd1 vccd1 _17320_/X sky130_fd_sc_hd__mux2_1
X_14532_ _15781_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14532_/Y sky130_fd_sc_hd__nor2_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26518_ _21122_/X _26518_/D vssd1 vssd1 vccd1 vccd1 _26518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27498_ _27726_/CLK _27498_/D vssd1 vssd1 vccd1 vccd1 _27498_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _26638_/Q _14460_/X _14455_/X _14462_/Y vssd1 vssd1 vccd1 vccd1 _26638_/D
+ sky130_fd_sc_hd__a31o_1
X_17251_ _17251_/A vssd1 vssd1 vccd1 vccd1 _27935_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26449_ _20884_/X _26449_/D vssd1 vssd1 vccd1 vccd1 _26449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13414_ _14804_/A vssd1 vssd1 vccd1 vccd1 _13414_/X sky130_fd_sc_hd__buf_4
X_16202_ _26049_/Q _16221_/B _16221_/C vssd1 vssd1 vccd1 vccd1 _16202_/X sky130_fd_sc_hd__and3_1
XFILLER_179_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17182_ _25825_/Q _26024_/Q _17219_/S vssd1 vssd1 vccd1 vccd1 _17182_/X sky130_fd_sc_hd__mux2_1
X_14394_ _14394_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14394_/Y sky130_fd_sc_hd__nor2_1
X_16133_ _27404_/Q _16298_/B vssd1 vssd1 vccd1 vccd1 _16133_/Y sky130_fd_sc_hd__nand2_1
X_13345_ _26994_/Q _13344_/X _13351_/S vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _16353_/A _16313_/B _16313_/C vssd1 vssd1 vccd1 vccd1 _16400_/A sky130_fd_sc_hd__nand3_2
XFILLER_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13276_ _27021_/Q _13128_/X _13280_/S vssd1 vssd1 vccd1 vccd1 _13277_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15015_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15015_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19823_ _19823_/A vssd1 vssd1 vccd1 vccd1 _19823_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19754_ _19745_/X _19747_/X _19749_/X _19751_/X _19752_/X _19753_/X vssd1 vssd1 vccd1
+ vccd1 _19755_/A sky130_fd_sc_hd__mux4_1
XFILLER_111_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16966_ _27608_/Q _24635_/A _16974_/A vssd1 vssd1 vccd1 vccd1 _16967_/C sky130_fd_sc_hd__a21o_1
X_18705_ _26015_/Q _17692_/X _18713_/S vssd1 vssd1 vccd1 vccd1 _18706_/A sky130_fd_sc_hd__mux2_1
X_15917_ _15918_/A vssd1 vssd1 vccd1 vccd1 _15917_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19685_ _19685_/A vssd1 vssd1 vccd1 vccd1 _19685_/X sky130_fd_sc_hd__clkbuf_1
X_16897_ _16902_/A _16600_/Y _16309_/Y vssd1 vssd1 vccd1 vccd1 _16897_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18636_ _18636_/A vssd1 vssd1 vccd1 vccd1 _25984_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15848_ _15848_/A vssd1 vssd1 vccd1 vccd1 _26077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18567_ _26969_/Q _26937_/Q _26905_/Q _26873_/Q _17841_/X _17843_/X vssd1 vssd1 vccd1
+ vccd1 _18567_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15779_ _15779_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15779_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _17517_/X _25840_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17519_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18498_ _18498_/A _18474_/X vssd1 vssd1 vccd1 vccd1 _18498_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17449_ _17449_/A vssd1 vssd1 vccd1 vccd1 _25818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20460_ _20445_/X _20447_/X _20449_/X _20451_/X _20452_/X _20453_/X vssd1 vssd1 vccd1
+ vccd1 _20461_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119_ _27804_/Q _26565_/Q _26437_/Q _26117_/Q _19118_/X _19019_/X vssd1 vssd1 vccd1
+ vccd1 _19119_/X sky130_fd_sc_hd__mux4_2
X_20391_ _20391_/A vssd1 vssd1 vccd1 vccd1 _20391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22130_ _22162_/A vssd1 vssd1 vccd1 vccd1 _22130_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22061_ _22051_/X _22052_/X _22053_/X _22054_/X _22055_/X _22056_/X vssd1 vssd1 vccd1
+ vccd1 _22062_/A sky130_fd_sc_hd__mux4_1
XFILLER_161_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21012_ _21028_/A vssd1 vssd1 vccd1 vccd1 _21012_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25820_ _25913_/CLK _25820_/D vssd1 vssd1 vccd1 vccd1 _25820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25751_ _17444_/X _27832_/Q _25757_/S vssd1 vssd1 vccd1 vccd1 _25752_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22963_ _22955_/X _22956_/X _22957_/X _22958_/X _22960_/X _22962_/X vssd1 vssd1 vccd1
+ vccd1 _22964_/A sky130_fd_sc_hd__mux4_1
XFILLER_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21914_ _21914_/A vssd1 vssd1 vccd1 vccd1 _21914_/X sky130_fd_sc_hd__clkbuf_1
X_24702_ _27182_/Q _24711_/B vssd1 vssd1 vccd1 vccd1 _24702_/X sky130_fd_sc_hd__or2_1
X_25682_ _25682_/A vssd1 vssd1 vccd1 vccd1 _25682_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22894_ _22958_/A vssd1 vssd1 vccd1 vccd1 _22894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24633_ _24633_/A _24636_/A _24633_/C vssd1 vssd1 vccd1 vccd1 _24634_/A sky130_fd_sc_hd__and3_1
XFILLER_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27421_ _27792_/CLK _27421_/D vssd1 vssd1 vccd1 vccd1 _27421_/Q sky130_fd_sc_hd__dfxtp_1
X_21845_ _22017_/A vssd1 vssd1 vccd1 vccd1 _21912_/A sky130_fd_sc_hd__buf_2
XFILLER_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24564_ _24564_/A vssd1 vssd1 vccd1 vccd1 _27543_/D sky130_fd_sc_hd__clkbuf_1
X_27352_ _27352_/CLK _27352_/D vssd1 vssd1 vccd1 vccd1 _27352_/Q sky130_fd_sc_hd__dfxtp_2
X_21776_ _21776_/A vssd1 vssd1 vccd1 vccd1 _21776_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26303_ _20373_/X _26303_/D vssd1 vssd1 vccd1 vccd1 _26303_/Q sky130_fd_sc_hd__dfxtp_1
X_23515_ _23515_/A vssd1 vssd1 vccd1 vccd1 _27196_/D sky130_fd_sc_hd__clkbuf_1
X_27283_ _27678_/CLK _27283_/D vssd1 vssd1 vccd1 vccd1 _27283_/Q sky130_fd_sc_hd__dfxtp_1
X_20727_ _20759_/A vssd1 vssd1 vccd1 vccd1 _20727_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24495_ _24631_/A _24495_/B vssd1 vssd1 vccd1 vccd1 _24496_/A sky130_fd_sc_hd__and2_1
XFILLER_168_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26234_ _20129_/X _26234_/D vssd1 vssd1 vccd1 vccd1 _26234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23446_ _27172_/Q _23456_/B vssd1 vssd1 vccd1 vccd1 _23446_/X sky130_fd_sc_hd__or2_1
XFILLER_184_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20658_ _20652_/X _20653_/X _20654_/X _20655_/X _20656_/X _20657_/X vssd1 vssd1 vccd1
+ vccd1 _20659_/A sky130_fd_sc_hd__mux4_1
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26165_ _19889_/X _26165_/D vssd1 vssd1 vccd1 vccd1 _26165_/Q sky130_fd_sc_hd__dfxtp_1
X_23377_ _27760_/Q vssd1 vssd1 vccd1 vccd1 _24752_/A sky130_fd_sc_hd__inv_2
XFILLER_99_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20589_ _20589_/A vssd1 vssd1 vccd1 vccd1 _20589_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25116_ _27690_/Q _25112_/X _25115_/Y _23498_/X vssd1 vssd1 vccd1 vccd1 _27690_/D
+ sky130_fd_sc_hd__o211a_1
X_13130_ _13130_/A vssd1 vssd1 vccd1 vccd1 _27053_/D sky130_fd_sc_hd__clkbuf_1
X_22328_ _22328_/A vssd1 vssd1 vccd1 vccd1 _22328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26096_ _19651_/X _26096_/D vssd1 vssd1 vccd1 vccd1 _26096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25047_ _27074_/Q _27106_/Q _25047_/S vssd1 vssd1 vccd1 vccd1 _25047_/X sky130_fd_sc_hd__mux2_1
X_13061_ _13061_/A vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__clkbuf_4
X_22259_ _22245_/X _22246_/X _22247_/X _22248_/X _22249_/X _22250_/X vssd1 vssd1 vccd1
+ vccd1 _22260_/A sky130_fd_sc_hd__mux4_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16820_ _16816_/Y _16819_/Y _16807_/Y vssd1 vssd1 vccd1 vccd1 _16820_/X sky130_fd_sc_hd__a21o_1
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26998_ _22798_/X _26998_/D vssd1 vssd1 vccd1 vccd1 _26998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16751_ _16751_/A _16751_/B vssd1 vssd1 vccd1 vccd1 _16751_/Y sky130_fd_sc_hd__nand2_1
X_13963_ _26805_/Q _13949_/X _13944_/X _13962_/Y vssd1 vssd1 vccd1 vccd1 _26805_/D
+ sky130_fd_sc_hd__a31o_1
X_25949_ _26051_/CLK _25949_/D vssd1 vssd1 vccd1 vccd1 _25949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15702_ _26136_/Q _15040_/X _15697_/X _15701_/Y vssd1 vssd1 vccd1 vccd1 _26136_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19470_ _19462_/X _19464_/X _19468_/X _19448_/X _19469_/X vssd1 vssd1 vccd1 vccd1
+ _19471_/C sky130_fd_sc_hd__a221o_1
X_13894_ _13920_/A vssd1 vssd1 vccd1 vccd1 _13904_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16682_ _16077_/A _16751_/A _16681_/B _16699_/A vssd1 vssd1 vccd1 vccd1 _16682_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18421_ _18419_/X _18420_/X _18488_/S vssd1 vssd1 vccd1 vccd1 _18421_/X sky130_fd_sc_hd__mux2_2
XFILLER_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27619_ _27700_/CLK _27619_/D vssd1 vssd1 vccd1 vccd1 _27619_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ _15633_/A vssd1 vssd1 vccd1 vccd1 _26166_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _18342_/X _18351_/X _18352_/S vssd1 vssd1 vccd1 vccd1 _18353_/B sky130_fd_sc_hd__mux2_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15621_/S vssd1 vssd1 vccd1 vccd1 _15573_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17303_/A vssd1 vssd1 vccd1 vccd1 _17303_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _14515_/A vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__clkbuf_2
X_18283_ _26411_/Q _26379_/Q _26347_/Q _26315_/Q _18189_/X _18214_/X vssd1 vssd1 vccd1
+ vccd1 _18283_/X sky130_fd_sc_hd__mux4_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _13094_/X _26227_/Q _15501_/S vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17234_ _27084_/Q _27116_/Q _17234_/S vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__mux2_1
X_14446_ _15718_/A _14446_/B vssd1 vssd1 vccd1 vccd1 _14446_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ _26664_/Q _14365_/X _14371_/X _14376_/Y vssd1 vssd1 vccd1 vccd1 _26664_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17165_ _17165_/A vssd1 vssd1 vccd1 vccd1 _27928_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_156_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16116_ _16252_/B vssd1 vssd1 vccd1 vccd1 _16274_/B sky130_fd_sc_hd__clkbuf_1
X_13328_ _14718_/A vssd1 vssd1 vccd1 vccd1 _13328_/X sky130_fd_sc_hd__buf_2
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17096_ _17094_/X _17096_/B vssd1 vssd1 vccd1 vccd1 _17096_/X sky130_fd_sc_hd__and2b_1
XFILLER_192_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16047_ _27474_/Q vssd1 vssd1 vccd1 vccd1 _16047_/Y sky130_fd_sc_hd__inv_2
X_13259_ _13259_/A vssd1 vssd1 vccd1 vccd1 _27029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19806_ _19796_/X _19797_/X _19798_/X _19799_/X _19800_/X _19801_/X vssd1 vssd1 vccd1
+ vccd1 _19807_/A sky130_fd_sc_hd__mux4_1
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17998_ _27799_/Q _26560_/Q _26432_/Q _26112_/Q _17996_/X _17997_/X vssd1 vssd1 vccd1
+ vccd1 _17998_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19737_ _19737_/A vssd1 vssd1 vccd1 vccd1 _19737_/X sky130_fd_sc_hd__clkbuf_1
X_16949_ _25430_/A _18584_/A _24828_/B vssd1 vssd1 vccd1 vccd1 _24511_/A sky130_fd_sc_hd__and3_4
XFILLER_38_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19668_ _19659_/X _19661_/X _19663_/X _19665_/X _19666_/X _19667_/X vssd1 vssd1 vccd1
+ vccd1 _19669_/A sky130_fd_sc_hd__mux4_1
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18619_ _18691_/A _23109_/A _25735_/B vssd1 vssd1 vccd1 vccd1 _18676_/A sky130_fd_sc_hd__and3b_1
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19599_ _19589_/X _19590_/X _19591_/X _19592_/X _19593_/X _19594_/X vssd1 vssd1 vccd1
+ vccd1 _19600_/A sky130_fd_sc_hd__mux4_1
X_21630_ _21630_/A vssd1 vssd1 vccd1 vccd1 _21630_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21561_ _21561_/A vssd1 vssd1 vccd1 vccd1 _21561_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23300_ _23300_/A _23300_/B _23299_/X vssd1 vssd1 vccd1 vccd1 _23309_/A sky130_fd_sc_hd__or3b_1
X_20512_ _20512_/A vssd1 vssd1 vccd1 vccd1 _20512_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24280_ _16228_/X _16229_/X _16230_/X _24279_/X vssd1 vssd1 vccd1 vccd1 _27416_/D
+ sky130_fd_sc_hd__o31a_1
X_21492_ _21492_/A vssd1 vssd1 vccd1 vccd1 _21492_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23231_ _17492_/X _27151_/Q _23237_/S vssd1 vssd1 vccd1 vccd1 _23232_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20443_ _20443_/A vssd1 vssd1 vccd1 vccd1 _20443_/X sky130_fd_sc_hd__clkbuf_1
X_23162_ _23162_/A vssd1 vssd1 vccd1 vccd1 _27120_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20374_ _20354_/X _20357_/X _20360_/X _20363_/X _20364_/X _20365_/X vssd1 vssd1 vccd1
+ vccd1 _20375_/A sky130_fd_sc_hd__mux4_1
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22113_ _22161_/A vssd1 vssd1 vccd1 vccd1 _22113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23093_ _23093_/A vssd1 vssd1 vccd1 vccd1 _27090_/D sky130_fd_sc_hd__clkbuf_1
X_27970_ _27970_/A _15951_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22044_ _22044_/A vssd1 vssd1 vccd1 vccd1 _22044_/X sky130_fd_sc_hd__clkbuf_1
X_26921_ _22530_/X _26921_/D vssd1 vssd1 vccd1 vccd1 _26921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26852_ _22294_/X _26852_/D vssd1 vssd1 vccd1 vccd1 _26852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25803_ _17520_/X _27856_/Q _25805_/S vssd1 vssd1 vccd1 vccd1 _25804_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23995_ _27787_/Q vssd1 vssd1 vccd1 vccd1 _24031_/S sky130_fd_sc_hd__clkbuf_2
X_26783_ _22048_/X _26783_/D vssd1 vssd1 vccd1 vccd1 _26783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22946_ _22946_/A vssd1 vssd1 vccd1 vccd1 _22946_/X sky130_fd_sc_hd__clkbuf_1
X_25734_ _25734_/A vssd1 vssd1 vccd1 vccd1 _27825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25665_ _25654_/X _25656_/X _25658_/X _25660_/X _25661_/X _25662_/X vssd1 vssd1 vccd1
+ vccd1 _25666_/A sky130_fd_sc_hd__mux4_1
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22877_ _22869_/X _22870_/X _22871_/X _22872_/X _22874_/X _22876_/X vssd1 vssd1 vccd1
+ vccd1 _22878_/A sky130_fd_sc_hd__mux4_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27404_ _27404_/CLK _27404_/D vssd1 vssd1 vccd1 vccd1 _27404_/Q sky130_fd_sc_hd__dfxtp_1
X_21828_ _21828_/A vssd1 vssd1 vccd1 vccd1 _21828_/X sky130_fd_sc_hd__clkbuf_1
X_24616_ _27667_/Q _24620_/B vssd1 vssd1 vccd1 vccd1 _24617_/A sky130_fd_sc_hd__and2_1
X_25596_ _27716_/Q _25433_/X _25435_/X vssd1 vssd1 vccd1 vccd1 _25596_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_169_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24547_ _24547_/A vssd1 vssd1 vccd1 vccd1 _27536_/D sky130_fd_sc_hd__clkbuf_1
X_27335_ _27335_/CLK _27335_/D vssd1 vssd1 vccd1 vccd1 _27335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21759_ _22017_/A vssd1 vssd1 vccd1 vccd1 _21826_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14300_ _14388_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14300_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15280_ _26322_/Q _13344_/X _15284_/S vssd1 vssd1 vccd1 vccd1 _15281_/A sky130_fd_sc_hd__mux2_1
X_24478_ _27636_/Q _24478_/B vssd1 vssd1 vccd1 vccd1 _24479_/A sky130_fd_sc_hd__and2_1
X_27266_ _27266_/CLK _27266_/D vssd1 vssd1 vccd1 vccd1 _27266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14231_ _26716_/Q _14225_/X _14220_/X _14230_/Y vssd1 vssd1 vccd1 vccd1 _26716_/D
+ sky130_fd_sc_hd__a31o_1
X_26217_ _20071_/X _26217_/D vssd1 vssd1 vccd1 vccd1 _26217_/Q sky130_fd_sc_hd__dfxtp_1
X_23429_ _23429_/A vssd1 vssd1 vccd1 vccd1 _23429_/X sky130_fd_sc_hd__buf_2
X_27197_ _27207_/CLK _27197_/D vssd1 vssd1 vccd1 vccd1 _27197_/Q sky130_fd_sc_hd__dfxtp_1
X_14162_ _14340_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14162_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26148_ _19827_/X _26148_/D vssd1 vssd1 vccd1 vccd1 _26148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _13113_/A vssd1 vssd1 vccd1 vccd1 _27056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14093_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14093_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18970_ _26687_/Q _26655_/Q _26623_/Q _26591_/Q _18847_/X _18939_/X vssd1 vssd1 vccd1
+ vccd1 _18970_/X sky130_fd_sc_hd__mux4_2
XFILLER_4_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26079_ _19588_/X _26079_/D vssd1 vssd1 vccd1 vccd1 _26079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _27796_/Q _26557_/Q _26429_/Q _26109_/Q _17920_/X _17785_/X vssd1 vssd1 vccd1
+ vccd1 _17921_/X sky130_fd_sc_hd__mux4_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _15334_/B _15045_/B _15334_/C vssd1 vssd1 vccd1 vccd1 _14885_/A sky130_fd_sc_hd__or3b_2
XFILLER_105_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17852_ _17844_/X _17849_/X _18568_/S vssd1 vssd1 vccd1 vccd1 _17852_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _16826_/A _16908_/B vssd1 vssd1 vccd1 vccd1 _16803_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_113_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17783_ _27594_/Q vssd1 vssd1 vccd1 vccd1 _18455_/A sky130_fd_sc_hd__clkbuf_2
X_14995_ _26445_/Q _14988_/X _14989_/X _14994_/Y vssd1 vssd1 vccd1 vccd1 _26445_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19522_ _19516_/X _19518_/X _19521_/X _18837_/X _19312_/S vssd1 vssd1 vccd1 vccd1
+ _19531_/B sky130_fd_sc_hd__a221o_1
X_16734_ _16733_/B _16734_/B vssd1 vssd1 vccd1 vccd1 _16734_/X sky130_fd_sc_hd__and2b_1
X_13946_ _13964_/A vssd1 vssd1 vccd1 vccd1 _13954_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19453_ _19534_/A _19453_/B vssd1 vssd1 vccd1 vccd1 _19453_/X sky130_fd_sc_hd__or2_1
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16665_ _16816_/A _16666_/B vssd1 vssd1 vccd1 vccd1 _16665_/X sky130_fd_sc_hd__and2_1
X_13877_ _26835_/Q _13865_/X _13873_/X _13876_/Y vssd1 vssd1 vccd1 vccd1 _26835_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_36 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18404_ _26961_/Q _26929_/Q _26897_/Q _26865_/Q _18403_/X _18269_/X vssd1 vssd1 vccd1
+ vccd1 _18404_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _15616_/A vssd1 vssd1 vccd1 vccd1 _26173_/D sky130_fd_sc_hd__clkbuf_1
X_19384_ _19409_/A _19384_/B vssd1 vssd1 vccd1 vccd1 _19384_/X sky130_fd_sc_hd__or2_1
X_16596_ _16835_/A _16596_/B vssd1 vssd1 vccd1 vccd1 _16599_/B sky130_fd_sc_hd__xnor2_1
XFILLER_201_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18335_ _26702_/Q _26670_/Q _26638_/Q _26606_/Q _18011_/A _18481_/A vssd1 vssd1 vccd1
+ vccd1 _18336_/A sky130_fd_sc_hd__mux4_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _13234_/X _26203_/Q _15549_/S vssd1 vssd1 vccd1 vccd1 _15548_/A sky130_fd_sc_hd__mux2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18266_ _18844_/A vssd1 vssd1 vccd1 vccd1 _18398_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_129_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15478_ _15478_/A vssd1 vssd1 vccd1 vccd1 _26234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17217_ _25929_/Q _25995_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17218_/B sky130_fd_sc_hd__mux2_1
X_14429_ _14436_/A vssd1 vssd1 vccd1 vccd1 _14504_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18197_ _18195_/X _18196_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18197_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17148_ _17120_/X _17147_/X _17098_/X vssd1 vssd1 vccd1 vccd1 _17148_/X sky130_fd_sc_hd__a21bo_1
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17079_ _27200_/Q _17077_/X _17128_/S vssd1 vssd1 vccd1 vccd1 _17080_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20090_ _20076_/X _20077_/X _20078_/X _20079_/X _20081_/X _20083_/X vssd1 vssd1 vccd1
+ vccd1 _20091_/A sky130_fd_sc_hd__mux4_1
XFILLER_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22800_ _22800_/A vssd1 vssd1 vccd1 vccd1 _22800_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23780_ _23778_/X _23779_/X _23795_/S vssd1 vssd1 vccd1 vccd1 _23780_/X sky130_fd_sc_hd__mux2_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20992_ _21040_/A vssd1 vssd1 vccd1 vccd1 _20992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22731_ _22716_/X _22718_/X _22720_/X _22722_/X _22723_/X _22724_/X vssd1 vssd1 vccd1
+ vccd1 _22732_/A sky130_fd_sc_hd__mux4_1
XFILLER_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25450_ _27692_/Q _25448_/X _25449_/X vssd1 vssd1 vccd1 vccd1 _25450_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_168_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22662_ _22662_/A vssd1 vssd1 vccd1 vccd1 _22662_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24401_ _24401_/A vssd1 vssd1 vccd1 vccd1 _27480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21613_ _21599_/X _21600_/X _21601_/X _21602_/X _21603_/X _21604_/X vssd1 vssd1 vccd1
+ vccd1 _21614_/A sky130_fd_sc_hd__mux4_1
X_25381_ _25381_/A vssd1 vssd1 vccd1 vccd1 _27730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_18 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22593_ _22609_/A vssd1 vssd1 vccd1 vccd1 _22593_/X sky130_fd_sc_hd__clkbuf_1
X_27120_ _27295_/CLK _27120_/D vssd1 vssd1 vccd1 vccd1 _27120_/Q sky130_fd_sc_hd__dfxtp_1
X_24332_ _24332_/A vssd1 vssd1 vccd1 vccd1 _27449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21544_ _21544_/A vssd1 vssd1 vccd1 vccd1 _21544_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27051_ _22986_/X _27051_/D vssd1 vssd1 vccd1 vccd1 _27051_/Q sky130_fd_sc_hd__dfxtp_1
X_24263_ _24263_/A _24264_/B vssd1 vssd1 vccd1 vccd1 _27405_/D sky130_fd_sc_hd__nor2_1
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21475_ _21475_/A vssd1 vssd1 vccd1 vccd1 _21475_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26002_ _26002_/CLK _26002_/D vssd1 vssd1 vccd1 vccd1 _26002_/Q sky130_fd_sc_hd__dfxtp_1
X_23214_ _23214_/A vssd1 vssd1 vccd1 vccd1 _27143_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20426_ _20426_/A vssd1 vssd1 vccd1 vccd1 _20426_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24194_ _24194_/A vssd1 vssd1 vccd1 vccd1 _27367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23145_ _23167_/A vssd1 vssd1 vccd1 vccd1 _23154_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20357_ _20425_/A vssd1 vssd1 vccd1 vccd1 _20357_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23076_ _23076_/A vssd1 vssd1 vccd1 vccd1 _27082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27953_ _27953_/A _15922_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
X_20288_ _20336_/A vssd1 vssd1 vccd1 vccd1 _20288_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22027_ _22016_/X _22018_/X _22020_/X _22022_/X _22023_/X _22024_/X vssd1 vssd1 vccd1
+ vccd1 _22028_/A sky130_fd_sc_hd__mux4_1
X_26904_ _22470_/X _26904_/D vssd1 vssd1 vccd1 vccd1 _26904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26835_ _22236_/X _26835_/D vssd1 vssd1 vccd1 vccd1 _26835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13800_ _26861_/Q _13793_/X _13794_/X _13799_/Y vssd1 vssd1 vccd1 vccd1 _26861_/D
+ sky130_fd_sc_hd__a31o_1
X_26766_ _21990_/X _26766_/D vssd1 vssd1 vccd1 vccd1 _26766_/Q sky130_fd_sc_hd__dfxtp_1
X_14780_ _14779_/X _26532_/Q _14789_/S vssd1 vssd1 vccd1 vccd1 _14781_/A sky130_fd_sc_hd__mux2_1
X_23978_ _23975_/X _23977_/X _23985_/S vssd1 vssd1 vccd1 vccd1 _23978_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13731_ _26886_/Q _13724_/X _13718_/X _13730_/Y vssd1 vssd1 vccd1 vccd1 _26886_/D
+ sky130_fd_sc_hd__a31o_1
X_25717_ _25705_/X _25706_/X _25707_/X _25708_/X _25709_/X _25710_/X vssd1 vssd1 vccd1
+ vccd1 _25718_/A sky130_fd_sc_hd__mux4_1
X_22929_ _22923_/X _22924_/X _22925_/X _22926_/X _22927_/X _22928_/X vssd1 vssd1 vccd1
+ vccd1 _22930_/A sky130_fd_sc_hd__mux4_1
X_26697_ _21752_/X _26697_/D vssd1 vssd1 vccd1 vccd1 _26697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16450_ _16450_/A _16450_/B vssd1 vssd1 vccd1 vccd1 _16450_/Y sky130_fd_sc_hd__xnor2_1
X_13662_ _26910_/Q _13653_/X _13656_/X _13661_/Y vssd1 vssd1 vccd1 vccd1 _26910_/D
+ sky130_fd_sc_hd__a31o_1
X_25648_ _25648_/A vssd1 vssd1 vccd1 vccd1 _25648_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _14804_/X _26268_/Q _15401_/S vssd1 vssd1 vccd1 vccd1 _15402_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _13861_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13593_/Y sky130_fd_sc_hd__nor2_1
X_16381_ _16751_/B _16398_/B vssd1 vssd1 vccd1 vccd1 _16383_/A sky130_fd_sc_hd__or2_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25579_ _27713_/Q _25568_/X _25569_/X vssd1 vssd1 vccd1 vccd1 _25579_/Y sky130_fd_sc_hd__a21oi_1
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18405_/A vssd1 vssd1 vccd1 vccd1 _18216_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_185_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15332_ _26298_/Q _13420_/X _15332_/S vssd1 vssd1 vccd1 vccd1 _15333_/A sky130_fd_sc_hd__mux2_1
X_27318_ _27323_/CLK _27318_/D vssd1 vssd1 vccd1 vccd1 _27318_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18051_ _18043_/X _18046_/X _18050_/X _18026_/X _17990_/X vssd1 vssd1 vccd1 vccd1
+ _18052_/C sky130_fd_sc_hd__a221o_1
X_27249_ _27264_/CLK _27249_/D vssd1 vssd1 vccd1 vccd1 _27249_/Q sky130_fd_sc_hd__dfxtp_1
X_15263_ _15319_/A vssd1 vssd1 vccd1 vccd1 _15332_/S sky130_fd_sc_hd__buf_2
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _16998_/X _17000_/X _17299_/A vssd1 vssd1 vccd1 vccd1 _17002_/X sky130_fd_sc_hd__a21bo_1
XFILLER_184_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14214_ _26723_/Q _14212_/X _14207_/X _14213_/Y vssd1 vssd1 vccd1 vccd1 _26723_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA_6 _21686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _15194_/A vssd1 vssd1 vccd1 vccd1 _26361_/D sky130_fd_sc_hd__clkbuf_1
X_14145_ _14410_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _14145_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14076_ _14090_/A vssd1 vssd1 vccd1 vccd1 _14076_/X sky130_fd_sc_hd__clkbuf_2
X_18953_ _27600_/Q vssd1 vssd1 vccd1 vccd1 _19485_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13027_ _13027_/A vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__clkbuf_2
X_17904_ _18000_/A vssd1 vssd1 vccd1 vccd1 _17904_/X sky130_fd_sc_hd__buf_6
X_18884_ _19004_/A _18884_/B vssd1 vssd1 vccd1 vccd1 _18884_/X sky130_fd_sc_hd__or2_1
XFILLER_94_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17835_ _18324_/A vssd1 vssd1 vccd1 vccd1 _17835_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17766_ _27436_/Q vssd1 vssd1 vccd1 vccd1 _17766_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14978_ _26452_/Q _14974_/X _14976_/X _14977_/Y vssd1 vssd1 vccd1 vccd1 _26452_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19505_ _26166_/Q _26102_/Q _27030_/Q _26998_/Q _19460_/X _19482_/X vssd1 vssd1 vccd1
+ vccd1 _19506_/B sky130_fd_sc_hd__mux4_1
X_16717_ _16731_/A _16731_/B _16433_/A vssd1 vssd1 vccd1 vccd1 _16719_/A sky130_fd_sc_hd__a21o_1
X_13929_ _26815_/Q _13919_/X _13925_/X _13928_/Y vssd1 vssd1 vccd1 vccd1 _26815_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17697_ _25918_/Q _17696_/X _17706_/S vssd1 vssd1 vccd1 vccd1 _17698_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19436_ _19434_/X _19435_/X _19480_/S vssd1 vssd1 vccd1 vccd1 _19436_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16648_ _16648_/A _16648_/B _16648_/C vssd1 vssd1 vccd1 vccd1 _16648_/X sky130_fd_sc_hd__and3_1
XFILLER_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19367_ _19365_/X _19366_/X _19499_/S vssd1 vssd1 vccd1 vccd1 _19367_/X sky130_fd_sc_hd__mux2_1
X_16579_ _27402_/Q _16312_/X _16314_/X _14727_/A vssd1 vssd1 vccd1 vccd1 _16579_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18318_ _18318_/A _18317_/X vssd1 vssd1 vccd1 vccd1 _18318_/X sky130_fd_sc_hd__or2b_1
XFILLER_175_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19298_ _26701_/Q _26669_/Q _26637_/Q _26605_/Q _19297_/X _19227_/A vssd1 vssd1 vccd1
+ vccd1 _19299_/B sky130_fd_sc_hd__mux4_2
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ _18408_/A vssd1 vssd1 vccd1 vccd1 _18249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_814 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21260_ _21260_/A vssd1 vssd1 vccd1 vccd1 _21260_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20211_ _20211_/A vssd1 vssd1 vccd1 vccd1 _20211_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21191_ _21179_/X _21180_/X _21181_/X _21182_/X _21183_/X _21184_/X vssd1 vssd1 vccd1
+ vccd1 _21192_/A sky130_fd_sc_hd__mux4_1
XFILLER_144_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27990__456 vssd1 vssd1 vccd1 vccd1 _27990__456/HI _27990_/A sky130_fd_sc_hd__conb_1
X_20142_ _20130_/X _20131_/X _20132_/X _20133_/X _20134_/X _20135_/X vssd1 vssd1 vccd1
+ vccd1 _20143_/A sky130_fd_sc_hd__mux4_1
XFILLER_44_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20073_ _20073_/A vssd1 vssd1 vccd1 vccd1 _20073_/X sky130_fd_sc_hd__clkbuf_1
X_24950_ _27666_/Q _24935_/X _24949_/Y _24938_/X vssd1 vssd1 vccd1 vccd1 _27666_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23901_ _27787_/Q vssd1 vssd1 vccd1 vccd1 _23938_/S sky130_fd_sc_hd__clkbuf_2
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24881_ _24877_/A _24880_/C _27766_/Q vssd1 vssd1 vccd1 vccd1 _24882_/B sky130_fd_sc_hd__a21oi_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater340 _27720_/CLK vssd1 vssd1 vccd1 vccd1 _27719_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26620_ _21484_/X _26620_/D vssd1 vssd1 vccd1 vccd1 _26620_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater351 _27582_/CLK vssd1 vssd1 vccd1 vccd1 _27754_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater362 _27576_/CLK vssd1 vssd1 vccd1 vccd1 _25909_/CLK sky130_fd_sc_hd__clkbuf_1
X_23832_ _27073_/Q _23812_/X _23813_/X _27105_/Q _23814_/X vssd1 vssd1 vccd1 vccd1
+ _23832_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater373 _27555_/CLK vssd1 vssd1 vccd1 vccd1 _27558_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater384 _27462_/CLK vssd1 vssd1 vccd1 vccd1 _27207_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater395 _27368_/CLK vssd1 vssd1 vccd1 vccd1 _27825_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23763_ _23861_/A vssd1 vssd1 vccd1 vccd1 _23763_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26551_ _21246_/X _26551_/D vssd1 vssd1 vccd1 vccd1 _26551_/Q sky130_fd_sc_hd__dfxtp_1
X_20975_ _21147_/A vssd1 vssd1 vccd1 vccd1 _21041_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25502_ _25500_/X _25199_/B _25501_/X _25483_/X vssd1 vssd1 vccd1 vccd1 _25502_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22714_ _22714_/A vssd1 vssd1 vccd1 vccd1 _22714_/X sky130_fd_sc_hd__clkbuf_1
X_23694_ _27772_/Q _27252_/Q _23694_/S vssd1 vssd1 vccd1 vccd1 _23695_/A sky130_fd_sc_hd__mux2_1
X_26482_ _21002_/X _26482_/D vssd1 vssd1 vccd1 vccd1 _26482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22645_ _22630_/X _22632_/X _22634_/X _22636_/X _22637_/X _22638_/X vssd1 vssd1 vccd1
+ vccd1 _22646_/A sky130_fd_sc_hd__mux4_1
X_25433_ _25539_/A vssd1 vssd1 vccd1 vccd1 _25433_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25364_ _25364_/A vssd1 vssd1 vccd1 vccd1 _27722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22576_ _22576_/A vssd1 vssd1 vccd1 vccd1 _22576_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27103_ _27103_/CLK _27103_/D vssd1 vssd1 vccd1 vccd1 _27103_/Q sky130_fd_sc_hd__dfxtp_1
X_21527_ _21513_/X _21514_/X _21515_/X _21516_/X _21517_/X _21518_/X vssd1 vssd1 vccd1
+ vccd1 _21528_/A sky130_fd_sc_hd__mux4_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24315_ _27542_/Q _24317_/B vssd1 vssd1 vccd1 vccd1 _24316_/A sky130_fd_sc_hd__and2_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25295_ _25295_/A _25295_/B vssd1 vssd1 vccd1 vccd1 _25296_/B sky130_fd_sc_hd__xnor2_1
XFILLER_181_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24246_ _24246_/A vssd1 vssd1 vccd1 vccd1 _27394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27034_ _22922_/X _27034_/D vssd1 vssd1 vccd1 vccd1 _27034_/Q sky130_fd_sc_hd__dfxtp_1
X_21458_ _21458_/A vssd1 vssd1 vccd1 vccd1 _21458_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20409_ _20425_/A vssd1 vssd1 vccd1 vccd1 _20409_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24177_ _24177_/A vssd1 vssd1 vccd1 vccd1 _27359_/D sky130_fd_sc_hd__clkbuf_1
X_21389_ _21389_/A vssd1 vssd1 vccd1 vccd1 _21389_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23128_ _27105_/Q _17699_/X _23132_/S vssd1 vssd1 vccd1 vccd1 _23129_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27936_ _27936_/A _15947_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
X_15950_ _15956_/A vssd1 vssd1 vccd1 vccd1 _15955_/A sky130_fd_sc_hd__buf_2
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23059_ _27075_/Q _17705_/X _23059_/S vssd1 vssd1 vccd1 vccd1 _23060_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14901_ _14731_/X _26483_/Q _14907_/S vssd1 vssd1 vccd1 vccd1 _14902_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ _15881_/A vssd1 vssd1 vccd1 vccd1 _15881_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17620_ _17620_/A vssd1 vssd1 vccd1 vccd1 _25882_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26818_ _22170_/X _26818_/D vssd1 vssd1 vccd1 vccd1 _26818_/Q sky130_fd_sc_hd__dfxtp_1
X_14832_ _14832_/A vssd1 vssd1 vccd1 vccd1 _26514_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27798_ _25646_/X _27798_/D vssd1 vssd1 vccd1 vccd1 _27798_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _17453_/X _25852_/Q _17551_/S vssd1 vssd1 vccd1 vccd1 _17552_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1094 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26749_ _21928_/X _26749_/D vssd1 vssd1 vccd1 vccd1 _26749_/Q sky130_fd_sc_hd__dfxtp_1
X_14763_ _16252_/A vssd1 vssd1 vccd1 vccd1 _14763_/X sky130_fd_sc_hd__buf_2
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _16502_/A _16508_/B vssd1 vssd1 vccd1 vccd1 _16502_/Y sky130_fd_sc_hd__nor2_1
X_13714_ _13895_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13714_/Y sky130_fd_sc_hd__nor2_1
X_17482_ _27426_/Q vssd1 vssd1 vccd1 vccd1 _17482_/X sky130_fd_sc_hd__clkbuf_2
X_14694_ _15767_/A _14699_/B vssd1 vssd1 vccd1 vccd1 _14694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19221_ _18801_/X _19215_/X _19217_/X _19219_/X _19220_/X vssd1 vssd1 vccd1 vccd1
+ _19222_/C sky130_fd_sc_hd__a221o_1
X_16433_ _16433_/A _16433_/B vssd1 vssd1 vccd1 vccd1 _16433_/Y sky130_fd_sc_hd__nor2_1
X_13645_ _13915_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19152_ _19143_/X _19146_/X _19150_/X _19151_/X _19105_/X vssd1 vssd1 vccd1 vccd1
+ _19153_/C sky130_fd_sc_hd__a221o_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _25949_/Q vssd1 vssd1 vccd1 vccd1 _16364_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ _14527_/A vssd1 vssd1 vccd1 vccd1 _13938_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _18437_/A vssd1 vssd1 vccd1 vccd1 _18197_/S sky130_fd_sc_hd__clkbuf_2
X_28004__470 vssd1 vssd1 vccd1 vccd1 _28004__470/HI _28004_/A sky130_fd_sc_hd__conb_1
X_15315_ _26306_/Q _13395_/X _15317_/S vssd1 vssd1 vccd1 vccd1 _15316_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19083_ _19107_/A _19083_/B _19083_/C vssd1 vssd1 vccd1 vccd1 _19084_/A sky130_fd_sc_hd__and3_1
X_16295_ _16151_/A _24305_/A _16845_/A vssd1 vssd1 vccd1 vccd1 _16583_/A sky130_fd_sc_hd__o21a_1
XFILLER_184_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18034_ _18085_/A vssd1 vssd1 vccd1 vccd1 _18034_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15246_ _15246_/A vssd1 vssd1 vccd1 vccd1 _26337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15177_ _15177_/A vssd1 vssd1 vccd1 vccd1 _26368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14128_ _14394_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_592 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19985_ _19985_/A vssd1 vssd1 vccd1 vccd1 _19985_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14059_ _14531_/A vssd1 vssd1 vccd1 vccd1 _14412_/A sky130_fd_sc_hd__clkbuf_2
X_18936_ _18936_/A vssd1 vssd1 vccd1 vccd1 _26045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18867_ _18858_/X _18861_/X _18865_/X _18866_/X _18840_/X vssd1 vssd1 vccd1 vccd1
+ _18868_/C sky130_fd_sc_hd__a221o_1
XFILLER_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17818_ _27597_/Q vssd1 vssd1 vccd1 vccd1 _18412_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18798_ _19492_/A vssd1 vssd1 vccd1 vccd1 _19560_/A sky130_fd_sc_hd__clkbuf_2
X_17749_ _17749_/A vssd1 vssd1 vccd1 vccd1 _25934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20760_ _20754_/X _20755_/X _20756_/X _20757_/X _20758_/X _20759_/X vssd1 vssd1 vccd1
+ vccd1 _20761_/A sky130_fd_sc_hd__mux4_1
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19419_ _19419_/A _19419_/B vssd1 vssd1 vccd1 vccd1 _19419_/X sky130_fd_sc_hd__or2_1
XFILLER_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20691_ _20759_/A vssd1 vssd1 vccd1 vccd1 _20691_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22430_ _22430_/A vssd1 vssd1 vccd1 vccd1 _22430_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22361_ _22347_/X _22348_/X _22349_/X _22350_/X _22352_/X _22354_/X vssd1 vssd1 vccd1
+ vccd1 _22362_/A sky130_fd_sc_hd__mux4_1
XFILLER_109_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24100_ _27398_/Q _24106_/B vssd1 vssd1 vccd1 vccd1 _24101_/A sky130_fd_sc_hd__and2_1
X_21312_ _21312_/A vssd1 vssd1 vccd1 vccd1 _21312_/X sky130_fd_sc_hd__clkbuf_1
X_25080_ _25078_/X _25079_/X _25087_/S vssd1 vssd1 vccd1 vccd1 _25080_/X sky130_fd_sc_hd__mux2_1
X_22292_ _22292_/A vssd1 vssd1 vccd1 vccd1 _22292_/X sky130_fd_sc_hd__clkbuf_1
X_24031_ _24029_/X _24030_/X _24031_/S vssd1 vssd1 vccd1 vccd1 _24031_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21243_ _21231_/X _21234_/X _21237_/X _21240_/X _21241_/X _21242_/X vssd1 vssd1 vccd1
+ vccd1 _21244_/A sky130_fd_sc_hd__mux4_1
XFILLER_151_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21174_ _21174_/A vssd1 vssd1 vccd1 vccd1 _21174_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20125_ _20125_/A vssd1 vssd1 vccd1 vccd1 _20125_/X sky130_fd_sc_hd__clkbuf_1
X_25982_ _27416_/CLK _25982_/D vssd1 vssd1 vccd1 vccd1 _25982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27721_ _27746_/CLK _27721_/D vssd1 vssd1 vccd1 vccd1 _27721_/Q sky130_fd_sc_hd__dfxtp_1
X_20056_ _20044_/X _20045_/X _20046_/X _20047_/X _20048_/X _20049_/X vssd1 vssd1 vccd1
+ vccd1 _20057_/A sky130_fd_sc_hd__mux4_1
X_24933_ _24937_/A _24933_/B vssd1 vssd1 vccd1 vccd1 _24933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27652_ _27654_/CLK _27652_/D vssd1 vssd1 vccd1 vccd1 _27652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24864_ _24914_/A vssd1 vssd1 vccd1 vccd1 _24864_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater170 _27112_/CLK vssd1 vssd1 vccd1 vccd1 _27081_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26603_ _21424_/X _26603_/D vssd1 vssd1 vccd1 vccd1 _26603_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater181 _27790_/CLK vssd1 vssd1 vccd1 vccd1 _27674_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _14500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23815_ _27071_/Q _23812_/X _23813_/X _27103_/Q _23814_/X vssd1 vssd1 vccd1 vccd1
+ _23815_/X sky130_fd_sc_hd__a221o_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater192 _25984_/CLK vssd1 vssd1 vccd1 vccd1 _27833_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27583_ _27584_/CLK _27583_/D vssd1 vssd1 vccd1 vccd1 _27583_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _14518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24795_ _27631_/Q _24785_/X _24794_/Y _24787_/X vssd1 vssd1 vccd1 vccd1 _27631_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _16756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _17356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26534_ _21178_/X _26534_/D vssd1 vssd1 vccd1 vccd1 _26534_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_248 _27773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 _26818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23746_ _27785_/Q vssd1 vssd1 vccd1 vccd1 _23946_/A sky130_fd_sc_hd__buf_2
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20958_ _21027_/A vssd1 vssd1 vccd1 vccd1 _20958_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26465_ _20944_/X _26465_/D vssd1 vssd1 vccd1 vccd1 _26465_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23677_ _27764_/Q _27244_/Q _23683_/S vssd1 vssd1 vccd1 vccd1 _23678_/A sky130_fd_sc_hd__mux2_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _21147_/A vssd1 vssd1 vccd1 vccd1 _20955_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25416_ _27746_/Q input58/X _25424_/S vssd1 vssd1 vccd1 vccd1 _25417_/A sky130_fd_sc_hd__mux2_1
X_13430_ _27366_/Q _13108_/A _13102_/A _27334_/Q _13036_/X vssd1 vssd1 vccd1 vccd1
+ _16033_/A sky130_fd_sc_hd__a221oi_4
XFILLER_167_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22628_ _22628_/A vssd1 vssd1 vccd1 vccd1 _22628_/X sky130_fd_sc_hd__clkbuf_1
X_26396_ _20695_/X _26396_/D vssd1 vssd1 vccd1 vccd1 _26396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13361_ _26989_/Q _13360_/X _13367_/S vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__mux2_1
X_22559_ _22539_/X _22542_/X _22545_/X _22548_/X _22549_/X _22550_/X vssd1 vssd1 vccd1
+ vccd1 _22560_/A sky130_fd_sc_hd__mux4_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25347_ _25347_/A _27517_/Q vssd1 vssd1 vccd1 vccd1 _25348_/B sky130_fd_sc_hd__or2_1
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15100_ _15100_/A vssd1 vssd1 vccd1 vccd1 _26402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16080_ _16559_/A _16845_/B _16073_/C vssd1 vssd1 vccd1 vccd1 _16602_/B sky130_fd_sc_hd__a21oi_1
X_13292_ _13292_/A vssd1 vssd1 vccd1 vccd1 _27014_/D sky130_fd_sc_hd__clkbuf_1
X_25278_ _25310_/A vssd1 vssd1 vccd1 vccd1 _25332_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15031_ _26432_/Q _15028_/X _15029_/X _15030_/Y vssd1 vssd1 vccd1 vccd1 _26432_/D
+ sky130_fd_sc_hd__a31o_1
X_27017_ _22864_/X _27017_/D vssd1 vssd1 vccd1 vccd1 _27017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24229_ _24229_/A vssd1 vssd1 vccd1 vccd1 _27384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19770_ _19764_/X _19765_/X _19766_/X _19767_/X _19768_/X _19769_/X vssd1 vssd1 vccd1
+ vccd1 _19771_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16982_ _16979_/A _24636_/A _16982_/C _16982_/D vssd1 vssd1 vccd1 vccd1 _16983_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18721_ _18721_/A vssd1 vssd1 vccd1 vccd1 _26022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27919_ _27919_/A _15970_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
X_15933_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15933_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18652_ _25992_/Q _17721_/X _18652_/S vssd1 vssd1 vccd1 vccd1 _18653_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _15868_/A vssd1 vssd1 vccd1 vccd1 _15864_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17603_ _17671_/S vssd1 vssd1 vccd1 vccd1 _17612_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _14883_/S vssd1 vssd1 vccd1 vccd1 _14824_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18583_ _18583_/A vssd1 vssd1 vccd1 vccd1 _25975_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _15795_/A vssd1 vssd1 vccd1 vccd1 _26101_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17534_ _17428_/X _25844_/Q _17540_/S vssd1 vssd1 vccd1 vccd1 _17535_/A sky130_fd_sc_hd__mux2_1
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14746_/A vssd1 vssd1 vccd1 vccd1 _26543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17465_ _17465_/A vssd1 vssd1 vccd1 vccd1 _25823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_199_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14677_ _15751_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14677_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19204_ _26825_/Q _26793_/Q _26761_/Q _26729_/Q _19203_/X _19111_/X vssd1 vssd1 vccd1
+ vccd1 _19205_/B sky130_fd_sc_hd__mux4_1
X_16416_ _16447_/B _16447_/C _16369_/X vssd1 vssd1 vccd1 vccd1 _16417_/B sky130_fd_sc_hd__o21a_1
X_13628_ _26923_/Q _13626_/X _13616_/X _13627_/Y vssd1 vssd1 vccd1 vccd1 _26923_/D
+ sky130_fd_sc_hd__a31o_1
X_17396_ _20796_/A vssd1 vssd1 vccd1 vccd1 _25657_/A sky130_fd_sc_hd__buf_6
X_19135_ _26694_/Q _26662_/Q _26630_/Q _26598_/Q _18908_/X _18909_/X vssd1 vssd1 vccd1
+ vccd1 _19136_/B sky130_fd_sc_hd__mux4_2
Xrepeater84 _27296_/CLK vssd1 vssd1 vccd1 vccd1 _27425_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater95 _25935_/CLK vssd1 vssd1 vccd1 vccd1 _26002_/CLK sky130_fd_sc_hd__clkbuf_1
X_16347_ _16862_/B _16347_/B vssd1 vssd1 vccd1 vccd1 _16347_/Y sky130_fd_sc_hd__nand2_1
X_13559_ _27340_/Q _13063_/A _13082_/X _27308_/Q _13208_/X vssd1 vssd1 vccd1 vccd1
+ _14515_/A sky130_fd_sc_hd__a221oi_4
XFILLER_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19066_ _19501_/A _19066_/B vssd1 vssd1 vccd1 vccd1 _19066_/X sky130_fd_sc_hd__or2_1
XFILLER_121_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16278_ _27537_/Q _16254_/S vssd1 vssd1 vccd1 vccd1 _16278_/X sky130_fd_sc_hd__or2b_1
XFILLER_173_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18017_ _17995_/X _18003_/X _18008_/X _18015_/X _18016_/X vssd1 vssd1 vccd1 vccd1
+ _18028_/B sky130_fd_sc_hd__a221o_1
XFILLER_145_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15229_ _15229_/A vssd1 vssd1 vccd1 vccd1 _26345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19968_ _19956_/X _19957_/X _19958_/X _19959_/X _19960_/X _19961_/X vssd1 vssd1 vccd1
+ vccd1 _19969_/A sky130_fd_sc_hd__mux4_1
XFILLER_68_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18919_ _18895_/X _18904_/X _18911_/X _18918_/X _18880_/X vssd1 vssd1 vccd1 vccd1
+ _18935_/B sky130_fd_sc_hd__a221o_1
XFILLER_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19899_ _19899_/A vssd1 vssd1 vccd1 vccd1 _19899_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21930_ _21997_/A vssd1 vssd1 vccd1 vccd1 _21930_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21861_ _21844_/X _21846_/X _21848_/X _21850_/X _21851_/X _21852_/X vssd1 vssd1 vccd1
+ vccd1 _21862_/A sky130_fd_sc_hd__mux4_1
XFILLER_36_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20812_ _20791_/X _20795_/X _20799_/X _20803_/X _20804_/X _20805_/X vssd1 vssd1 vccd1
+ vccd1 _20813_/A sky130_fd_sc_hd__mux4_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23600_ _23600_/A vssd1 vssd1 vccd1 vccd1 _23616_/S sky130_fd_sc_hd__clkbuf_2
X_21792_ _21792_/A vssd1 vssd1 vccd1 vccd1 _21792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24580_ _24580_/A vssd1 vssd1 vccd1 vccd1 _27550_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20743_ _20759_/A vssd1 vssd1 vccd1 vccd1 _20743_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23531_ _23543_/A _23531_/B vssd1 vssd1 vccd1 vccd1 _23532_/A sky130_fd_sc_hd__and2_1
XFILLER_168_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26250_ _20191_/X _26250_/D vssd1 vssd1 vccd1 vccd1 _26250_/Q sky130_fd_sc_hd__dfxtp_1
X_23462_ input15/X _23455_/X _23459_/X _23461_/X vssd1 vssd1 vccd1 vccd1 _27177_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20674_ _20668_/X _20669_/X _20670_/X _20671_/X _20672_/X _20673_/X vssd1 vssd1 vccd1
+ vccd1 _20675_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22413_ _22401_/X _22402_/X _22403_/X _22404_/X _22405_/X _22406_/X vssd1 vssd1 vccd1
+ vccd1 _22414_/A sky130_fd_sc_hd__mux4_1
X_25201_ _27531_/Q _27499_/Q vssd1 vssd1 vccd1 vccd1 _25203_/A sky130_fd_sc_hd__nand2_1
XFILLER_183_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23393_ _23393_/A _23393_/B _23393_/C _23393_/D vssd1 vssd1 vccd1 vccd1 _23410_/C
+ sky130_fd_sc_hd__or4_1
X_26181_ _19949_/X _26181_/D vssd1 vssd1 vccd1 vccd1 _26181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22344_ _22344_/A vssd1 vssd1 vccd1 vccd1 _22344_/X sky130_fd_sc_hd__clkbuf_1
X_25132_ _25132_/A vssd1 vssd1 vccd1 vccd1 _25132_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27996__462 vssd1 vssd1 vccd1 vccd1 _27996__462/HI _27996_/A sky130_fd_sc_hd__conb_1
XFILLER_191_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25063_ _25922_/Q _25988_/Q _25821_/Q _26020_/Q _25052_/X _25027_/X vssd1 vssd1 vccd1
+ vccd1 _25063_/X sky130_fd_sc_hd__mux4_1
X_22275_ _22261_/X _22262_/X _22263_/X _22264_/X _22266_/X _22268_/X vssd1 vssd1 vccd1
+ vccd1 _22276_/A sky130_fd_sc_hd__mux4_1
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24014_ _24014_/A vssd1 vssd1 vccd1 vccd1 _24014_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21226_ _21226_/A vssd1 vssd1 vccd1 vccd1 _21226_/X sky130_fd_sc_hd__clkbuf_1
X_21157_ _21144_/X _21146_/X _21148_/X _21150_/X _21151_/X _21152_/X vssd1 vssd1 vccd1
+ vccd1 _21158_/A sky130_fd_sc_hd__mux4_1
XFILLER_137_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20108_ _20095_/X _20097_/X _20099_/X _20101_/X _20102_/X _20103_/X vssd1 vssd1 vccd1
+ vccd1 _20109_/A sky130_fd_sc_hd__mux4_1
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21088_ _21088_/A vssd1 vssd1 vccd1 vccd1 _21088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25965_ _26053_/CLK _25965_/D vssd1 vssd1 vccd1 vccd1 _25965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27704_ _27705_/CLK _27704_/D vssd1 vssd1 vccd1 vccd1 _27704_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24916_ _24940_/A vssd1 vssd1 vccd1 vccd1 _24937_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_20039_ _20039_/A vssd1 vssd1 vccd1 vccd1 _20039_/X sky130_fd_sc_hd__clkbuf_1
X_12930_ input9/X _27859_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _12931_/B sky130_fd_sc_hd__mux2_1
X_25896_ _25897_/CLK _25896_/D vssd1 vssd1 vccd1 vccd1 _25896_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27635_ _27636_/CLK _27635_/D vssd1 vssd1 vccd1 vccd1 _27635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24847_ _27645_/Q _24834_/X _24846_/Y _24839_/X vssd1 vssd1 vccd1 vccd1 _27645_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _15762_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14600_/Y sky130_fd_sc_hd__nor2_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _26189_/Q _14750_/A _15584_/S vssd1 vssd1 vccd1 vccd1 _15581_/A sky130_fd_sc_hd__mux2_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27566_ _27569_/CLK _27566_/D vssd1 vssd1 vccd1 vccd1 _27566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24778_ _24778_/A _24786_/B vssd1 vssd1 vccd1 vccd1 _24778_/Y sky130_fd_sc_hd__nand2_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14531_ _14531_/A vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__buf_2
XFILLER_18_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26517_ _21120_/X _26517_/D vssd1 vssd1 vccd1 vccd1 _26517_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23729_ _24063_/A vssd1 vssd1 vccd1 vccd1 _24050_/B sky130_fd_sc_hd__clkbuf_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27497_ _27726_/CLK _27497_/D vssd1 vssd1 vccd1 vccd1 _27497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17250_ _27214_/Q _17249_/X _17250_/S vssd1 vssd1 vccd1 vccd1 _17251_/A sky130_fd_sc_hd__mux2_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _15730_/A _14465_/B vssd1 vssd1 vccd1 vccd1 _14462_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26448_ _20882_/X _26448_/D vssd1 vssd1 vccd1 vccd1 _26448_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16201_ _16201_/A vssd1 vssd1 vccd1 vccd1 _16221_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_139_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13413_ _13413_/A vssd1 vssd1 vccd1 vccd1 _26973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17181_ _17181_/A vssd1 vssd1 vccd1 vccd1 _17181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14393_ _14393_/A vssd1 vssd1 vccd1 vccd1 _14403_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_26379_ _20635_/X _26379_/D vssd1 vssd1 vccd1 vccd1 _26379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16132_ _16132_/A vssd1 vssd1 vccd1 vccd1 _16298_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13344_ _14734_/A vssd1 vssd1 vccd1 vccd1 _13344_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _16057_/X _16063_/B _16063_/C _16063_/D vssd1 vssd1 vccd1 vccd1 _16313_/C
+ sky130_fd_sc_hd__and4b_1
X_13275_ _13275_/A vssd1 vssd1 vccd1 vccd1 _27022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_560 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15014_ _26438_/Q _15002_/X _15003_/X _15013_/Y vssd1 vssd1 vccd1 vccd1 _26438_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19822_ _19812_/X _19813_/X _19814_/X _19815_/X _19817_/X _19819_/X vssd1 vssd1 vccd1
+ vccd1 _19823_/A sky130_fd_sc_hd__mux4_1
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19753_ _19801_/A vssd1 vssd1 vccd1 vccd1 _19753_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16965_ _27592_/Q _27591_/Q _27590_/Q _16960_/A vssd1 vssd1 vccd1 vccd1 _16974_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_110_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _18761_/S vssd1 vssd1 vccd1 vccd1 _18713_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15916_ _15918_/A vssd1 vssd1 vccd1 vccd1 _15916_/Y sky130_fd_sc_hd__inv_2
X_19684_ _19678_/X _19679_/X _19680_/X _19681_/X _19682_/X _19683_/X vssd1 vssd1 vccd1
+ vccd1 _19685_/A sky130_fd_sc_hd__mux4_1
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16896_ _24240_/A _16896_/B _16896_/C _16895_/X vssd1 vssd1 vccd1 vccd1 _25582_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18635_ _25984_/Q _17696_/X _18641_/S vssd1 vssd1 vccd1 vccd1 _18636_/A sky130_fd_sc_hd__mux2_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _13222_/X _26077_/Q _15849_/S vssd1 vssd1 vccd1 vccd1 _15848_/A sky130_fd_sc_hd__mux2_1
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18566_ _27824_/Q _26585_/Q _26457_/Q _26137_/Q _17789_/X _17791_/X vssd1 vssd1 vccd1
+ vccd1 _18566_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _26108_/Q _15774_/X _15766_/X _15777_/Y vssd1 vssd1 vccd1 vccd1 _26108_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17517_ _27437_/Q vssd1 vssd1 vccd1 vccd1 _17517_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14729_ _14727_/X _26548_/Q _14741_/S vssd1 vssd1 vccd1 vccd1 _14730_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18497_ _26709_/Q _26677_/Q _26645_/Q _26613_/Q _18345_/X _18408_/X vssd1 vssd1 vccd1
+ vccd1 _18498_/A sky130_fd_sc_hd__mux4_1
X_17448_ _17447_/X _25818_/Q _17454_/S vssd1 vssd1 vccd1 vccd1 _17449_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17379_ _27857_/Q _27161_/Q _25906_/Q _25874_/Q _17061_/A _17181_/A vssd1 vssd1 vccd1
+ vccd1 _17379_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19118_ _19465_/A vssd1 vssd1 vccd1 vccd1 _19118_/X sky130_fd_sc_hd__buf_2
XFILLER_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20390_ _20376_/X _20377_/X _20378_/X _20379_/X _20380_/X _20381_/X vssd1 vssd1 vccd1
+ vccd1 _20391_/A sky130_fd_sc_hd__mux4_1
XFILLER_146_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19049_ _19165_/A vssd1 vssd1 vccd1 vccd1 _19049_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22060_ _22060_/A vssd1 vssd1 vccd1 vccd1 _22060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21011_ _21027_/A vssd1 vssd1 vccd1 vccd1 _21011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25750_ _25750_/A vssd1 vssd1 vccd1 vccd1 _27831_/D sky130_fd_sc_hd__clkbuf_1
X_22962_ _23030_/A vssd1 vssd1 vccd1 vccd1 _22962_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24701_ _25434_/A vssd1 vssd1 vccd1 vccd1 _24711_/B sky130_fd_sc_hd__clkbuf_1
X_21913_ _21913_/A vssd1 vssd1 vccd1 vccd1 _21913_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25681_ _25673_/X _25674_/X _25675_/X _25676_/X _25677_/X _25678_/X vssd1 vssd1 vccd1
+ vccd1 _25682_/A sky130_fd_sc_hd__mux4_1
XFILLER_71_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22893_ _22893_/A vssd1 vssd1 vccd1 vccd1 _22958_/A sky130_fd_sc_hd__buf_2
X_27420_ _27420_/CLK _27420_/D vssd1 vssd1 vccd1 vccd1 _27420_/Q sky130_fd_sc_hd__dfxtp_1
X_24632_ _24632_/A vssd1 vssd1 vccd1 vccd1 _27574_/D sky130_fd_sc_hd__clkbuf_1
X_21844_ _21911_/A vssd1 vssd1 vccd1 vccd1 _21844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27351_ _27353_/CLK _27351_/D vssd1 vssd1 vccd1 vccd1 _27351_/Q sky130_fd_sc_hd__dfxtp_2
X_21775_ _21758_/X _21760_/X _21762_/X _21764_/X _21765_/X _21766_/X vssd1 vssd1 vccd1
+ vccd1 _21776_/A sky130_fd_sc_hd__mux4_1
X_24563_ _27643_/Q _24565_/B vssd1 vssd1 vccd1 vccd1 _24564_/A sky130_fd_sc_hd__and2_1
X_26302_ _20371_/X _26302_/D vssd1 vssd1 vccd1 vccd1 _26302_/Q sky130_fd_sc_hd__dfxtp_1
X_20726_ _20758_/A vssd1 vssd1 vccd1 vccd1 _20726_/X sky130_fd_sc_hd__clkbuf_2
X_23514_ _23526_/A _23514_/B vssd1 vssd1 vccd1 vccd1 _23515_/A sky130_fd_sc_hd__and2_1
XFILLER_168_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27282_ _27788_/CLK _27282_/D vssd1 vssd1 vccd1 vccd1 _27282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24494_ _24398_/A _24505_/B _24492_/Y _24629_/B _27585_/Q vssd1 vssd1 vccd1 vccd1
+ _24495_/B sky130_fd_sc_hd__a32o_1
X_26233_ _20127_/X _26233_/D vssd1 vssd1 vccd1 vccd1 _26233_/Q sky130_fd_sc_hd__dfxtp_1
X_23445_ _23500_/B vssd1 vssd1 vccd1 vccd1 _23456_/B sky130_fd_sc_hd__clkbuf_1
X_20657_ _20673_/A vssd1 vssd1 vccd1 vccd1 _20657_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23376_ _27236_/Q vssd1 vssd1 vccd1 vccd1 _23376_/Y sky130_fd_sc_hd__inv_2
X_26164_ _19881_/X _26164_/D vssd1 vssd1 vccd1 vccd1 _26164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20588_ _20582_/X _20583_/X _20584_/X _20585_/X _20586_/X _20587_/X vssd1 vssd1 vccd1
+ vccd1 _20589_/A sky130_fd_sc_hd__mux4_2
XFILLER_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25115_ _25115_/A _25356_/A vssd1 vssd1 vccd1 vccd1 _25115_/Y sky130_fd_sc_hd__nand2_1
X_22327_ _22315_/X _22316_/X _22317_/X _22318_/X _22319_/X _22320_/X vssd1 vssd1 vccd1
+ vccd1 _22328_/A sky130_fd_sc_hd__mux4_1
XFILLER_178_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26095_ _19649_/X _26095_/D vssd1 vssd1 vccd1 vccd1 _26095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ _13060_/A vssd1 vssd1 vccd1 vccd1 _27064_/D sky130_fd_sc_hd__clkbuf_1
X_22258_ _22258_/A vssd1 vssd1 vccd1 vccd1 _22258_/X sky130_fd_sc_hd__clkbuf_1
X_25046_ _25044_/X _25045_/X _25046_/S vssd1 vssd1 vccd1 vccd1 _25046_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21209_ _21195_/X _21196_/X _21197_/X _21198_/X _21199_/X _21200_/X vssd1 vssd1 vccd1
+ vccd1 _21210_/A sky130_fd_sc_hd__mux4_1
XFILLER_78_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22189_ _22173_/X _22174_/X _22175_/X _22176_/X _22179_/X _22182_/X vssd1 vssd1 vccd1
+ vccd1 _22190_/A sky130_fd_sc_hd__mux4_1
XFILLER_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26997_ _22796_/X _26997_/D vssd1 vssd1 vccd1 vccd1 _26997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16750_ _16743_/Y _16748_/X _16765_/D vssd1 vssd1 vccd1 vccd1 _16750_/X sky130_fd_sc_hd__a21o_1
X_13962_ _14342_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _13962_/Y sky130_fd_sc_hd__nor2_1
X_25948_ _26049_/CLK _25948_/D vssd1 vssd1 vccd1 vccd1 _25948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15701_ _15701_/A _15703_/B vssd1 vssd1 vccd1 vccd1 _15701_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16681_ _16751_/A _16681_/B vssd1 vssd1 vccd1 vccd1 _16681_/X sky130_fd_sc_hd__or2_1
XFILLER_100_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13893_ _13919_/A vssd1 vssd1 vccd1 vccd1 _13893_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25879_ _27383_/CLK _25879_/D vssd1 vssd1 vccd1 vccd1 _25879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18420_ _26417_/Q _26385_/Q _26353_/Q _26321_/Q _18305_/X _18329_/X vssd1 vssd1 vccd1
+ vccd1 _18420_/X sky130_fd_sc_hd__mux4_1
X_27618_ _27621_/CLK _27618_/D vssd1 vssd1 vccd1 vccd1 _27618_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _13072_/X _26166_/Q _15634_/S vssd1 vssd1 vccd1 vccd1 _15633_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18344_/X _18347_/X _18350_/X _18468_/A vssd1 vssd1 vccd1 vccd1 _18351_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27549_ _27659_/CLK _27549_/D vssd1 vssd1 vccd1 vccd1 _27549_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15563_/A vssd1 vssd1 vccd1 vccd1 _26197_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17277_/X _17302_/B vssd1 vssd1 vccd1 vccd1 _17302_/X sky130_fd_sc_hd__and2b_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14514_ _14530_/A vssd1 vssd1 vccd1 vccd1 _14514_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _26539_/Q _26507_/Q _26475_/Q _27051_/Q _18233_/X _18259_/X vssd1 vssd1 vccd1
+ vccd1 _18282_/X sky130_fd_sc_hd__mux4_1
XFILLER_70_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15494_/A vssd1 vssd1 vccd1 vccd1 _26228_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17233_ _17177_/X _17227_/X _17229_/X _17232_/X vssd1 vssd1 vccd1 vccd1 _17233_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14445_ _16563_/A vssd1 vssd1 vccd1 vccd1 _15718_/A sky130_fd_sc_hd__buf_2
XFILLER_30_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17164_ _27207_/Q _17163_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17165_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ _14376_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14376_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16115_ _16235_/B vssd1 vssd1 vccd1 vccd1 _16252_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13327_ _13327_/A vssd1 vssd1 vccd1 vccd1 _27000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17095_ _25919_/Q _25985_/Q _17132_/S vssd1 vssd1 vccd1 vccd1 _17096_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16046_ _16043_/Y _16044_/X _16045_/X vssd1 vssd1 vccd1 vccd1 _16066_/B sky130_fd_sc_hd__a21oi_1
X_13258_ _27029_/Q _13078_/X _13258_/S vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13189_ _16230_/A vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__buf_2
XFILLER_9_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19805_ _19805_/A vssd1 vssd1 vccd1 vccd1 _19805_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17997_ _18486_/A vssd1 vssd1 vccd1 vccd1 _17997_/X sky130_fd_sc_hd__buf_2
XFILLER_81_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19736_ _19726_/X _19727_/X _19728_/X _19729_/X _19731_/X _19733_/X vssd1 vssd1 vccd1
+ vccd1 _19737_/A sky130_fd_sc_hd__mux4_1
X_16948_ _25358_/A _24640_/A vssd1 vssd1 vccd1 vccd1 _24828_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ _16879_/A _16879_/B _16879_/C vssd1 vssd1 vccd1 vccd1 _16879_/X sky130_fd_sc_hd__and3_1
XFILLER_53_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19667_ _19715_/A vssd1 vssd1 vccd1 vccd1 _19667_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18618_ _18589_/X _18615_/X _18617_/Y _18604_/Y vssd1 vssd1 vccd1 vccd1 _25977_/D
+ sky130_fd_sc_hd__o211a_1
X_19598_ _19598_/A vssd1 vssd1 vccd1 vccd1 _19598_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18549_ _26968_/Q _26936_/Q _26904_/Q _26872_/Q _17841_/X _18427_/X vssd1 vssd1 vccd1
+ vccd1 _18549_/X sky130_fd_sc_hd__mux4_1
XFILLER_127_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21560_ _21560_/A vssd1 vssd1 vccd1 vccd1 _21560_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20511_ _20511_/A vssd1 vssd1 vccd1 vccd1 _20511_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21491_ _21475_/X _21476_/X _21477_/X _21478_/X _21480_/X _21482_/X vssd1 vssd1 vccd1
+ vccd1 _21492_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23230_ _23230_/A vssd1 vssd1 vccd1 vccd1 _27150_/D sky130_fd_sc_hd__clkbuf_1
X_20442_ _20424_/X _20425_/X _20426_/X _20427_/X _20430_/X _20433_/X vssd1 vssd1 vccd1
+ vccd1 _20443_/A sky130_fd_sc_hd__mux4_1
XFILLER_146_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23161_ _27120_/Q _17747_/X _23165_/S vssd1 vssd1 vccd1 vccd1 _23162_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20373_ _20373_/A vssd1 vssd1 vccd1 vccd1 _20373_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22112_ _22176_/A vssd1 vssd1 vccd1 vccd1 _22112_/X sky130_fd_sc_hd__clkbuf_1
X_23092_ _27090_/Q _17753_/X _23092_/S vssd1 vssd1 vccd1 vccd1 _23093_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22043_ _22035_/X _22036_/X _22037_/X _22038_/X _22039_/X _22040_/X vssd1 vssd1 vccd1
+ vccd1 _22044_/A sky130_fd_sc_hd__mux4_1
X_26920_ _22528_/X _26920_/D vssd1 vssd1 vccd1 vccd1 _26920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26851_ _22292_/X _26851_/D vssd1 vssd1 vccd1 vccd1 _26851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25802_ _25802_/A vssd1 vssd1 vccd1 vccd1 _27855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26782_ _22046_/X _26782_/D vssd1 vssd1 vccd1 vccd1 _26782_/Q sky130_fd_sc_hd__dfxtp_1
X_23994_ _25937_/Q _26003_/Q _25836_/Q _26035_/Q _23993_/X _23976_/X vssd1 vssd1 vccd1
+ vccd1 _23994_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25733_ _25733_/A _25733_/B vssd1 vssd1 vccd1 vccd1 _25734_/A sky130_fd_sc_hd__and2_1
X_22945_ _22939_/X _22940_/X _22941_/X _22942_/X _22943_/X _22944_/X vssd1 vssd1 vccd1
+ vccd1 _22946_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25664_ _25664_/A vssd1 vssd1 vccd1 vccd1 _25664_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22876_ _22944_/A vssd1 vssd1 vccd1 vccd1 _22876_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27403_ _27406_/CLK _27403_/D vssd1 vssd1 vccd1 vccd1 _27403_/Q sky130_fd_sc_hd__dfxtp_1
X_24615_ _24615_/A vssd1 vssd1 vccd1 vccd1 _27566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21827_ _21827_/A vssd1 vssd1 vccd1 vccd1 _21827_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25595_ _18594_/A _25326_/B _25594_/X _25566_/X vssd1 vssd1 vccd1 vccd1 _25595_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27334_ _27334_/CLK _27334_/D vssd1 vssd1 vccd1 vccd1 _27334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24546_ _24552_/A _24546_/B vssd1 vssd1 vccd1 vccd1 _24547_/A sky130_fd_sc_hd__and2_1
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21758_ _21825_/A vssd1 vssd1 vccd1 vccd1 _21758_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20709_ _20773_/A vssd1 vssd1 vccd1 vccd1 _20709_/X sky130_fd_sc_hd__clkbuf_1
X_27265_ _27266_/CLK _27265_/D vssd1 vssd1 vccd1 vccd1 _27265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24477_ _24477_/A vssd1 vssd1 vccd1 vccd1 _27514_/D sky130_fd_sc_hd__clkbuf_1
X_21689_ _21737_/A vssd1 vssd1 vccd1 vccd1 _21689_/X sky130_fd_sc_hd__clkbuf_1
X_14230_ _14408_/A _14234_/B vssd1 vssd1 vccd1 vccd1 _14230_/Y sky130_fd_sc_hd__nor2_1
X_26216_ _20069_/X _26216_/D vssd1 vssd1 vccd1 vccd1 _26216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23428_ input34/X _23415_/X _23427_/X _23421_/X vssd1 vssd1 vccd1 vccd1 _27165_/D
+ sky130_fd_sc_hd__o211a_1
X_27196_ _27196_/CLK _27196_/D vssd1 vssd1 vccd1 vccd1 _27196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14161_ _14215_/A vssd1 vssd1 vccd1 vccd1 _14174_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26147_ _19825_/X _26147_/D vssd1 vssd1 vccd1 vccd1 _26147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23359_ _24925_/A _23354_/Y _27261_/Q _24808_/A _23358_/X vssd1 vssd1 vccd1 vccd1
+ _23360_/C sky130_fd_sc_hd__o221a_1
XFILLER_153_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13112_ _27056_/Q _13111_/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ _26768_/Q _14090_/X _14080_/X _14091_/Y vssd1 vssd1 vccd1 vccd1 _26768_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26078_ _19586_/X _26078_/D vssd1 vssd1 vccd1 vccd1 _26078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17920_ _18401_/A vssd1 vssd1 vccd1 vccd1 _17920_/X sky130_fd_sc_hd__clkbuf_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _27270_/Q vssd1 vssd1 vccd1 vccd1 _15334_/C sky130_fd_sc_hd__buf_2
X_25029_ _25026_/X _25028_/X _25046_/S vssd1 vssd1 vccd1 vccd1 _25029_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17851_ _18405_/A vssd1 vssd1 vccd1 vccd1 _18568_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_132_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16802_ _16802_/A _16822_/A vssd1 vssd1 vccd1 vccd1 _16802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17782_ _18458_/A vssd1 vssd1 vccd1 vccd1 _17782_/X sky130_fd_sc_hd__buf_4
X_14994_ _15732_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14994_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19521_ _19519_/X _19520_/X _19539_/S vssd1 vssd1 vccd1 vccd1 _19521_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16733_ _16734_/B _16733_/B vssd1 vssd1 vccd1 vccd1 _16733_/X sky130_fd_sc_hd__and2b_1
X_13945_ _16033_/A vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19452_ _26836_/Q _26804_/Q _26772_/Q _26740_/Q _19338_/X _19407_/X vssd1 vssd1 vccd1
+ vccd1 _19453_/B sky130_fd_sc_hd__mux4_1
X_16664_ _16664_/A _16664_/B vssd1 vssd1 vccd1 vccd1 _16664_/X sky130_fd_sc_hd__xor2_1
X_13876_ _13876_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18403_ _18403_/A vssd1 vssd1 vccd1 vccd1 _18403_/X sky130_fd_sc_hd__clkbuf_2
X_15615_ _26173_/Q _14801_/A _15617_/S vssd1 vssd1 vccd1 vccd1 _15616_/A sky130_fd_sc_hd__mux2_1
X_19383_ _26833_/Q _26801_/Q _26769_/Q _26737_/Q _19338_/X _19248_/X vssd1 vssd1 vccd1
+ vccd1 _19384_/B sky130_fd_sc_hd__mux4_2
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16595_ _16639_/A _16595_/B vssd1 vssd1 vccd1 vccd1 _16596_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _18334_/A vssd1 vssd1 vccd1 vccd1 _25963_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15546_ _15546_/A vssd1 vssd1 vccd1 vccd1 _26204_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18265_ _18265_/A vssd1 vssd1 vccd1 vccd1 _25960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15477_ _26234_/Q _13420_/X _15477_/S vssd1 vssd1 vccd1 vccd1 _15478_/A sky130_fd_sc_hd__mux2_1
X_17216_ _17338_/A vssd1 vssd1 vccd1 vccd1 _17216_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14428_ _16134_/A vssd1 vssd1 vccd1 vccd1 _15708_/A sky130_fd_sc_hd__buf_2
XFILLER_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18196_ _26952_/Q _26920_/Q _26888_/Q _26856_/Q _18101_/X _18129_/X vssd1 vssd1 vccd1
+ vccd1 _18196_/X sky130_fd_sc_hd__mux4_2
XFILLER_190_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17147_ _25822_/Q _26021_/Q _17158_/S vssd1 vssd1 vccd1 vccd1 _17147_/X sky130_fd_sc_hd__mux2_1
X_14359_ _14359_/A _14363_/B vssd1 vssd1 vccd1 vccd1 _14359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17078_ _17387_/S vssd1 vssd1 vccd1 vccd1 _17128_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16029_ _27407_/Q _16144_/B vssd1 vssd1 vccd1 vccd1 _16029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19719_ _19719_/A vssd1 vssd1 vccd1 vccd1 _19719_/X sky130_fd_sc_hd__clkbuf_1
X_20991_ _21039_/A vssd1 vssd1 vccd1 vccd1 _20991_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22730_ _22730_/A vssd1 vssd1 vccd1 vccd1 _22730_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22661_ _22649_/X _22650_/X _22651_/X _22652_/X _22653_/X _22654_/X vssd1 vssd1 vccd1
+ vccd1 _22662_/A sky130_fd_sc_hd__mux4_1
XFILLER_129_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24400_ _24400_/A _24400_/B vssd1 vssd1 vccd1 vccd1 _24401_/A sky130_fd_sc_hd__and2_1
X_21612_ _21612_/A vssd1 vssd1 vccd1 vccd1 _21612_/X sky130_fd_sc_hd__clkbuf_1
X_25380_ _27730_/Q input72/X _25380_/S vssd1 vssd1 vccd1 vccd1 _25381_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22592_ _22592_/A vssd1 vssd1 vccd1 vccd1 _22592_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24331_ _27549_/Q _24339_/B vssd1 vssd1 vccd1 vccd1 _24332_/A sky130_fd_sc_hd__and2_1
X_21543_ _21529_/X _21530_/X _21531_/X _21532_/X _21533_/X _21534_/X vssd1 vssd1 vccd1
+ vccd1 _21544_/A sky130_fd_sc_hd__mux4_1
XFILLER_193_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27050_ _22984_/X _27050_/D vssd1 vssd1 vccd1 vccd1 _27050_/Q sky130_fd_sc_hd__dfxtp_1
X_21474_ _21474_/A vssd1 vssd1 vccd1 vccd1 _21474_/X sky130_fd_sc_hd__clkbuf_1
X_24262_ _24262_/A _24264_/B vssd1 vssd1 vccd1 vccd1 _27404_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_28021__487 vssd1 vssd1 vccd1 vccd1 _28021__487/HI _28021_/A sky130_fd_sc_hd__conb_1
X_26001_ _26001_/CLK _26001_/D vssd1 vssd1 vccd1 vccd1 _26001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23213_ _17466_/X _27143_/Q _23215_/S vssd1 vssd1 vccd1 vccd1 _23214_/A sky130_fd_sc_hd__mux2_1
X_20425_ _20425_/A vssd1 vssd1 vccd1 vccd1 _20425_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24193_ _27472_/Q _24195_/B vssd1 vssd1 vccd1 vccd1 _24194_/A sky130_fd_sc_hd__and2_1
XFILLER_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23144_ _23144_/A vssd1 vssd1 vccd1 vccd1 _27112_/D sky130_fd_sc_hd__clkbuf_1
X_20356_ _20704_/A vssd1 vssd1 vccd1 vccd1 _20425_/A sky130_fd_sc_hd__buf_2
XFILLER_49_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27952_ _27952_/A _15923_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
X_23075_ _27082_/Q _17728_/X _23081_/S vssd1 vssd1 vccd1 vccd1 _23076_/A sky130_fd_sc_hd__mux2_1
X_20287_ _20335_/A vssd1 vssd1 vccd1 vccd1 _20287_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22026_ _22026_/A vssd1 vssd1 vccd1 vccd1 _22026_/X sky130_fd_sc_hd__clkbuf_1
X_26903_ _22468_/X _26903_/D vssd1 vssd1 vccd1 vccd1 _26903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26834_ _22228_/X _26834_/D vssd1 vssd1 vccd1 vccd1 _26834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26765_ _21988_/X _26765_/D vssd1 vssd1 vccd1 vccd1 _26765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23977_ _25935_/Q _26001_/Q _25834_/Q _26033_/Q _23946_/X _23976_/X vssd1 vssd1 vccd1
+ vccd1 _23977_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _13910_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13730_/Y sky130_fd_sc_hd__nor2_1
X_25716_ _25716_/A vssd1 vssd1 vccd1 vccd1 _25716_/X sky130_fd_sc_hd__clkbuf_1
X_22928_ _22944_/A vssd1 vssd1 vccd1 vccd1 _22928_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26696_ _21750_/X _26696_/D vssd1 vssd1 vccd1 vccd1 _26696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _13930_/A _13661_/B vssd1 vssd1 vccd1 vccd1 _13661_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25647_ _25635_/X _25636_/X _25637_/X _25638_/X _25640_/X _25642_/X vssd1 vssd1 vccd1
+ vccd1 _25648_/A sky130_fd_sc_hd__mux4_1
X_22859_ _22853_/X _22854_/X _22855_/X _22856_/X _22857_/X _22858_/X vssd1 vssd1 vccd1
+ vccd1 _22860_/A sky130_fd_sc_hd__mux4_1
X_15400_ _15400_/A vssd1 vssd1 vccd1 vccd1 _26269_/D sky130_fd_sc_hd__clkbuf_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _16751_/A _16380_/B vssd1 vssd1 vccd1 vccd1 _16398_/B sky130_fd_sc_hd__xor2_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _26936_/Q _13580_/X _13587_/X _13591_/Y vssd1 vssd1 vccd1 vccd1 _26936_/D
+ sky130_fd_sc_hd__a31o_1
X_25578_ _18594_/X _25306_/B _25577_/X _18591_/X vssd1 vssd1 vccd1 vccd1 _25578_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _15331_/A vssd1 vssd1 vccd1 vccd1 _26299_/D sky130_fd_sc_hd__clkbuf_1
X_27317_ _27323_/CLK _27317_/D vssd1 vssd1 vccd1 vccd1 _27317_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24529_ _24529_/A vssd1 vssd1 vccd1 vccd1 _27531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18050_ _18047_/X _18049_/X _18075_/S vssd1 vssd1 vccd1 vccd1 _18050_/X sky130_fd_sc_hd__mux2_2
XFILLER_177_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27248_ _27250_/CLK _27248_/D vssd1 vssd1 vccd1 vccd1 _27248_/Q sky130_fd_sc_hd__dfxtp_1
X_15262_ _15551_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15319_/A sky130_fd_sc_hd__nor2_4
XFILLER_32_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17001_ input37/X vssd1 vssd1 vccd1 vccd1 _17299_/A sky130_fd_sc_hd__buf_2
XFILLER_172_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14213_ _14390_/A _14213_/B vssd1 vssd1 vccd1 vccd1 _14213_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27179_ _27180_/CLK _27179_/D vssd1 vssd1 vccd1 vccd1 _27179_/Q sky130_fd_sc_hd__dfxtp_1
X_15193_ _14709_/X _26361_/Q _15201_/S vssd1 vssd1 vccd1 vccd1 _15194_/A sky130_fd_sc_hd__mux2_1
XANTENNA_7 _21698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14144_ _26748_/Q _14142_/X _14133_/X _14143_/Y vssd1 vssd1 vccd1 vccd1 _26748_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14075_ _26774_/Q _14058_/X _14064_/X _14074_/Y vssd1 vssd1 vccd1 vccd1 _26774_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18952_ _19004_/A _18952_/B vssd1 vssd1 vccd1 vccd1 _18952_/X sky130_fd_sc_hd__or2_1
XFILLER_106_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17903_ _18462_/A vssd1 vssd1 vccd1 vccd1 _17903_/X sky130_fd_sc_hd__buf_6
X_13026_ _13081_/A vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__buf_2
XFILLER_105_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18883_ _26140_/Q _26076_/Q _27004_/Q _26972_/Q _18882_/X _18810_/X vssd1 vssd1 vccd1
+ vccd1 _18884_/B sky130_fd_sc_hd__mux4_1
XFILLER_117_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17834_ _18408_/A vssd1 vssd1 vccd1 vccd1 _18324_/A sky130_fd_sc_hd__buf_2
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17765_ _17765_/A vssd1 vssd1 vccd1 vccd1 _25939_/D sky130_fd_sc_hd__clkbuf_1
X_14977_ _15714_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19504_ _18895_/X _19499_/X _19501_/X _19503_/X _19312_/S vssd1 vssd1 vccd1 vccd1
+ _19513_/B sky130_fd_sc_hd__a221o_1
X_13928_ _13928_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _13928_/Y sky130_fd_sc_hd__nor2_1
X_16716_ _16383_/A _16393_/Y _16397_/X _16398_/X vssd1 vssd1 vccd1 vccd1 _16731_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17696_ _27414_/Q vssd1 vssd1 vccd1 vccd1 _17696_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19435_ _27818_/Q _26579_/Q _26451_/Q _26131_/Q _19414_/X _19321_/X vssd1 vssd1 vccd1
+ vccd1 _19435_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16647_ _16647_/A vssd1 vssd1 vccd1 vccd1 _16647_/X sky130_fd_sc_hd__buf_2
X_13859_ _13859_/A _13861_/B vssd1 vssd1 vccd1 vccd1 _13859_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16578_ _16916_/A _16585_/B vssd1 vssd1 vccd1 vccd1 _16578_/Y sky130_fd_sc_hd__nor2_1
X_19366_ _27815_/Q _26576_/Q _26448_/Q _26128_/Q _18922_/X _18901_/X vssd1 vssd1 vccd1
+ vccd1 _19366_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18317_ _18474_/A vssd1 vssd1 vccd1 vccd1 _18317_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15529_ _15529_/A vssd1 vssd1 vccd1 vccd1 _26212_/D sky130_fd_sc_hd__clkbuf_1
X_19297_ _19297_/A vssd1 vssd1 vccd1 vccd1 _19297_/X sky130_fd_sc_hd__buf_6
XFILLER_148_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _26826_/Q _26794_/Q _26762_/Q _26730_/Q _18175_/X _18199_/X vssd1 vssd1 vccd1
+ vccd1 _18248_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_826 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ _18179_/A _18156_/X vssd1 vssd1 vccd1 vccd1 _18179_/X sky130_fd_sc_hd__or2b_1
XFILLER_163_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20210_ _20200_/X _20201_/X _20202_/X _20203_/X _20204_/X _20205_/X vssd1 vssd1 vccd1
+ vccd1 _20211_/A sky130_fd_sc_hd__mux4_1
X_21190_ _21190_/A vssd1 vssd1 vccd1 vccd1 _21190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20141_ _20141_/A vssd1 vssd1 vccd1 vccd1 _20141_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20072_ _20060_/X _20061_/X _20062_/X _20063_/X _20064_/X _20065_/X vssd1 vssd1 vccd1
+ vccd1 _20073_/A sky130_fd_sc_hd__mux4_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23900_ _25927_/Q _25993_/Q _25826_/Q _26025_/Q _23899_/X _23882_/X vssd1 vssd1 vccd1
+ vccd1 _23900_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24880_ _27766_/Q _27765_/Q _24880_/C vssd1 vssd1 vccd1 vccd1 _24887_/B sky130_fd_sc_hd__and3_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater330 _27716_/CLK vssd1 vssd1 vccd1 vccd1 _27773_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater341 _27758_/CLK vssd1 vssd1 vccd1 vccd1 _27720_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater352 _27577_/CLK vssd1 vssd1 vccd1 vccd1 _27582_/CLK sky130_fd_sc_hd__clkbuf_1
X_23831_ _23829_/X _23830_/X _23846_/S vssd1 vssd1 vccd1 vccd1 _23831_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater363 _27681_/CLK vssd1 vssd1 vccd1 vccd1 _27379_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater374 _27651_/CLK vssd1 vssd1 vccd1 vccd1 _27555_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater385 _27105_/CLK vssd1 vssd1 vccd1 vccd1 _27350_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater396 _27473_/CLK vssd1 vssd1 vccd1 vccd1 _27368_/CLK sky130_fd_sc_hd__clkbuf_1
X_26550_ _21244_/X _26550_/D vssd1 vssd1 vccd1 vccd1 _26550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23762_ _24002_/A vssd1 vssd1 vccd1 vccd1 _23861_/A sky130_fd_sc_hd__buf_2
XFILLER_122_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ _21040_/A vssd1 vssd1 vccd1 vccd1 _20974_/X sky130_fd_sc_hd__clkbuf_1
X_25501_ _25487_/X _25492_/X _25493_/X _24875_/B _25494_/X vssd1 vssd1 vccd1 vccd1
+ _25501_/X sky130_fd_sc_hd__o311a_1
XFILLER_54_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22713_ _22697_/X _22698_/X _22699_/X _22700_/X _22702_/X _22704_/X vssd1 vssd1 vccd1
+ vccd1 _22714_/A sky130_fd_sc_hd__mux4_1
X_26481_ _21000_/X _26481_/D vssd1 vssd1 vccd1 vccd1 _26481_/Q sky130_fd_sc_hd__dfxtp_1
X_23693_ _23693_/A vssd1 vssd1 vccd1 vccd1 _27251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25432_ _27688_/Q vssd1 vssd1 vccd1 vccd1 _25539_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22644_ _22644_/A vssd1 vssd1 vccd1 vccd1 _22644_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25363_ _27722_/Q input52/X _25369_/S vssd1 vssd1 vccd1 vccd1 _25364_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22575_ _22561_/X _22562_/X _22563_/X _22564_/X _22565_/X _22566_/X vssd1 vssd1 vccd1
+ vccd1 _22576_/A sky130_fd_sc_hd__mux4_1
XFILLER_55_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27102_ _27413_/CLK _27102_/D vssd1 vssd1 vccd1 vccd1 _27102_/Q sky130_fd_sc_hd__dfxtp_1
X_24314_ _24314_/A vssd1 vssd1 vccd1 vccd1 _27441_/D sky130_fd_sc_hd__clkbuf_1
X_21526_ _21526_/A vssd1 vssd1 vccd1 vccd1 _21526_/X sky130_fd_sc_hd__clkbuf_1
X_25294_ _25299_/A _25290_/B _25287_/B vssd1 vssd1 vccd1 vccd1 _25295_/B sky130_fd_sc_hd__o21ai_1
XFILLER_194_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27033_ _22920_/X _27033_/D vssd1 vssd1 vccd1 vccd1 _27033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24245_ _24245_/A _24250_/B vssd1 vssd1 vccd1 vccd1 _24246_/A sky130_fd_sc_hd__and2_1
XFILLER_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21457_ _21443_/X _21444_/X _21445_/X _21446_/X _21447_/X _21448_/X vssd1 vssd1 vccd1
+ vccd1 _21458_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20408_ _20424_/A vssd1 vssd1 vccd1 vccd1 _20408_/X sky130_fd_sc_hd__clkbuf_1
X_21388_ _21388_/A vssd1 vssd1 vccd1 vccd1 _21388_/X sky130_fd_sc_hd__clkbuf_1
X_24176_ _27464_/Q _24184_/B vssd1 vssd1 vccd1 vccd1 _24177_/A sky130_fd_sc_hd__and2_1
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23127_ _23127_/A vssd1 vssd1 vccd1 vccd1 _27104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20339_ _20412_/A vssd1 vssd1 vccd1 vccd1 _20339_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27935_ _27935_/A _15948_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
X_23058_ _23058_/A vssd1 vssd1 vccd1 vccd1 _27074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_788 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14900_ _14900_/A vssd1 vssd1 vccd1 vccd1 _26484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22009_ _21997_/X _21998_/X _21999_/X _22000_/X _22002_/X _22004_/X vssd1 vssd1 vccd1
+ vccd1 _22010_/A sky130_fd_sc_hd__mux4_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _15881_/A vssd1 vssd1 vccd1 vccd1 _15880_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _26514_/Q _13344_/X _14835_/S vssd1 vssd1 vccd1 vccd1 _14832_/A sky130_fd_sc_hd__mux2_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26817_ _22168_/X _26817_/D vssd1 vssd1 vccd1 vccd1 _26817_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27797_ _25644_/X _27797_/D vssd1 vssd1 vccd1 vccd1 _27797_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17550_ _17550_/A vssd1 vssd1 vccd1 vccd1 _25851_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26748_ _21926_/X _26748_/D vssd1 vssd1 vccd1 vccd1 _26748_/Q sky130_fd_sc_hd__dfxtp_1
X_14762_ _14762_/A vssd1 vssd1 vccd1 vccd1 _26538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16501_ _16501_/A vssd1 vssd1 vccd1 vccd1 _16501_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13740_/A vssd1 vssd1 vccd1 vccd1 _13725_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17481_ _17481_/A vssd1 vssd1 vccd1 vccd1 _25828_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26679_ _21688_/X _26679_/D vssd1 vssd1 vccd1 vccd1 _26679_/Q sky130_fd_sc_hd__dfxtp_1
X_14693_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14693_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19220_ _19220_/A vssd1 vssd1 vccd1 vccd1 _19220_/X sky130_fd_sc_hd__clkbuf_2
X_16432_ _16890_/B _16719_/C vssd1 vssd1 vccd1 vccd1 _16433_/B sky130_fd_sc_hd__or2_1
X_13644_ _26917_/Q _13639_/X _13642_/X _13643_/Y vssd1 vssd1 vccd1 vccd1 _26917_/D
+ sky130_fd_sc_hd__a31o_1
X_19151_ _19290_/A vssd1 vssd1 vccd1 vccd1 _19151_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16395_/A _16395_/B vssd1 vssd1 vccd1 vccd1 _16851_/B sky130_fd_sc_hd__nor2_1
X_13575_ _27336_/Q _13108_/X _13029_/A _27304_/Q _13231_/X vssd1 vssd1 vccd1 vccd1
+ _14527_/A sky130_fd_sc_hd__a221oi_4
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ _26948_/Q _26916_/Q _26884_/Q _26852_/Q _18101_/X _17951_/X vssd1 vssd1 vccd1
+ vccd1 _18102_/X sky130_fd_sc_hd__mux4_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A vssd1 vssd1 vccd1 vccd1 _26307_/D sky130_fd_sc_hd__clkbuf_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ _19072_/X _19077_/X _19081_/X _19035_/X _18987_/X vssd1 vssd1 vccd1 vccd1
+ _19083_/C sky130_fd_sc_hd__a221o_1
XFILLER_157_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16294_ _26068_/Q _16137_/X _16293_/X vssd1 vssd1 vccd1 vccd1 _24305_/A sky130_fd_sc_hd__a21oi_2
XFILLER_173_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18033_ _18031_/X _18032_/X _18056_/S vssd1 vssd1 vccd1 vccd1 _18033_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _14788_/X _26337_/Q _15245_/S vssd1 vssd1 vccd1 vccd1 _15246_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15176_ _26368_/Q _13401_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15177_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _14127_/A vssd1 vssd1 vccd1 vccd1 _14138_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19984_ _19972_/X _19973_/X _19974_/X _19975_/X _19976_/X _19977_/X vssd1 vssd1 vccd1
+ vccd1 _19985_/A sky130_fd_sc_hd__mux4_1
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14058_ _14090_/A vssd1 vssd1 vccd1 vccd1 _14058_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18935_ _18989_/A _18935_/B _18935_/C vssd1 vssd1 vccd1 vccd1 _18936_/A sky130_fd_sc_hd__and3_1
XFILLER_122_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13009_ _27794_/Q _13009_/B vssd1 vssd1 vccd1 vccd1 _13010_/A sky130_fd_sc_hd__and2_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18866_ _19290_/A vssd1 vssd1 vccd1 vccd1 _18866_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17817_ _17799_/X _17806_/X _17814_/X _24394_/A vssd1 vssd1 vccd1 vccd1 _17817_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18797_ _18945_/A vssd1 vssd1 vccd1 vccd1 _19492_/A sky130_fd_sc_hd__clkbuf_4
X_17748_ _25934_/Q _17747_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17749_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17679_ _17679_/A vssd1 vssd1 vccd1 vccd1 _25912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1159 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19418_ _26162_/Q _26098_/Q _27026_/Q _26994_/Q _19326_/X _19348_/X vssd1 vssd1 vccd1
+ vccd1 _19419_/B sky130_fd_sc_hd__mux4_1
X_20690_ _20776_/A vssd1 vssd1 vccd1 vccd1 _20759_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19349_ _26159_/Q _26095_/Q _27023_/Q _26991_/Q _19326_/X _19348_/X vssd1 vssd1 vccd1
+ vccd1 _19350_/B sky130_fd_sc_hd__mux4_1
XFILLER_148_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22360_ _22360_/A vssd1 vssd1 vccd1 vccd1 _22360_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21311_ _21301_/X _21302_/X _21303_/X _21304_/X _21307_/X _21310_/X vssd1 vssd1 vccd1
+ vccd1 _21312_/A sky130_fd_sc_hd__mux4_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22291_ _22280_/X _22282_/X _22284_/X _22286_/X _22287_/X _22288_/X vssd1 vssd1 vccd1
+ vccd1 _22292_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24030_ _25941_/Q _26007_/Q _25840_/Q _26039_/Q _23993_/X _23744_/A vssd1 vssd1 vccd1
+ vccd1 _24030_/X sky130_fd_sc_hd__mux4_1
X_21242_ _21290_/A vssd1 vssd1 vccd1 vccd1 _21242_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21173_ _21163_/X _21164_/X _21165_/X _21166_/X _21167_/X _21168_/X vssd1 vssd1 vccd1
+ vccd1 _21174_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20124_ _20114_/X _20115_/X _20116_/X _20117_/X _20118_/X _20119_/X vssd1 vssd1 vccd1
+ vccd1 _20125_/A sky130_fd_sc_hd__mux4_1
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25981_ _26014_/CLK _25981_/D vssd1 vssd1 vccd1 vccd1 _25981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27720_ _27720_/CLK _27720_/D vssd1 vssd1 vccd1 vccd1 _27720_/Q sky130_fd_sc_hd__dfxtp_1
X_20055_ _20055_/A vssd1 vssd1 vccd1 vccd1 _20055_/X sky130_fd_sc_hd__clkbuf_1
X_24932_ _24941_/C _24932_/B vssd1 vssd1 vccd1 vccd1 _24933_/B sky130_fd_sc_hd__or2_1
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27651_ _27651_/CLK _27651_/D vssd1 vssd1 vccd1 vccd1 _27651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24863_ _24863_/A _24863_/B vssd1 vssd1 vccd1 vccd1 _24863_/Y sky130_fd_sc_hd__nand2_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_515 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater160 _27133_/CLK vssd1 vssd1 vccd1 vccd1 _27830_/CLK sky130_fd_sc_hd__clkbuf_1
X_26602_ _21422_/X _26602_/D vssd1 vssd1 vccd1 vccd1 _26602_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater171 _27111_/CLK vssd1 vssd1 vccd1 vccd1 _27112_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23814_ _23862_/A vssd1 vssd1 vccd1 vccd1 _23814_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater182 _27415_/CLK vssd1 vssd1 vccd1 vccd1 _27413_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27582_ _27582_/CLK _27582_/D vssd1 vssd1 vccd1 vccd1 _27582_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _14503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24794_ _24794_/A _24800_/B vssd1 vssd1 vccd1 vccd1 _24794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater193 _25985_/CLK vssd1 vssd1 vccd1 vccd1 _25984_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_199_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_216 _14524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 _25582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26533_ _21176_/X _26533_/D vssd1 vssd1 vccd1 vccd1 _26533_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23745_ _27826_/Q _27130_/Q _25875_/Q _25843_/Q _23997_/A _23744_/X vssd1 vssd1 vccd1
+ vccd1 _23745_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _17356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_249 _27773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ _21215_/A vssd1 vssd1 vccd1 vccd1 _21027_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26464_ _20936_/X _26464_/D vssd1 vssd1 vccd1 vccd1 _26464_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23676_ _23676_/A vssd1 vssd1 vccd1 vccd1 _27243_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20888_ _20954_/A vssd1 vssd1 vccd1 vccd1 _20888_/X sky130_fd_sc_hd__clkbuf_1
X_25415_ _25415_/A vssd1 vssd1 vccd1 vccd1 _25424_/S sky130_fd_sc_hd__buf_2
XFILLER_198_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22627_ _22609_/X _22610_/X _22611_/X _22612_/X _22615_/X _22618_/X vssd1 vssd1 vccd1
+ vccd1 _22628_/A sky130_fd_sc_hd__mux4_1
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26395_ _20693_/X _26395_/D vssd1 vssd1 vccd1 vccd1 _26395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25346_ _25354_/A _27517_/Q vssd1 vssd1 vccd1 vccd1 _25348_/A sky130_fd_sc_hd__nand2_1
X_13360_ _14750_/A vssd1 vssd1 vccd1 vccd1 _13360_/X sky130_fd_sc_hd__buf_2
XFILLER_195_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22558_ _22558_/A vssd1 vssd1 vccd1 vccd1 _22558_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21509_ _21494_/X _21496_/X _21498_/X _21500_/X _21501_/X _21502_/X vssd1 vssd1 vccd1
+ vccd1 _21510_/A sky130_fd_sc_hd__mux4_1
X_25277_ _27539_/Q vssd1 vssd1 vccd1 vccd1 _25310_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13291_ _27014_/Q _13166_/X _13291_/S vssd1 vssd1 vccd1 vccd1 _13292_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22489_ _22521_/A vssd1 vssd1 vccd1 vccd1 _22489_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15030_ _15767_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15030_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27016_ _22862_/X _27016_/D vssd1 vssd1 vccd1 vccd1 _27016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24228_ _24228_/A _24233_/B vssd1 vssd1 vccd1 vccd1 _24229_/A sky130_fd_sc_hd__and2_1
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24159_ _24159_/A vssd1 vssd1 vccd1 vccd1 _27351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16981_ _16981_/A vssd1 vssd1 vccd1 vccd1 _25909_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18720_ _26022_/Q _17715_/X _18724_/S vssd1 vssd1 vccd1 vccd1 _18721_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27918_ _27918_/A _15971_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15932_ _15956_/A vssd1 vssd1 vccd1 vccd1 _15937_/A sky130_fd_sc_hd__buf_2
XFILLER_114_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18651_ _18651_/A vssd1 vssd1 vccd1 vccd1 _25991_/D sky130_fd_sc_hd__clkbuf_1
X_15863_ _15988_/A vssd1 vssd1 vccd1 vccd1 _15868_/A sky130_fd_sc_hd__buf_4
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27849_ _27849_/CLK _27849_/D vssd1 vssd1 vccd1 vccd1 _27849_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _17658_/A vssd1 vssd1 vccd1 vccd1 _17671_/S sky130_fd_sc_hd__buf_2
X_14814_ _14870_/A vssd1 vssd1 vccd1 vccd1 _14883_/S sky130_fd_sc_hd__buf_2
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15794_ _13078_/X _26101_/Q _15794_/S vssd1 vssd1 vccd1 vccd1 _15795_/A sky130_fd_sc_hd__mux2_1
X_18582_ _18842_/A _18582_/B _18582_/C vssd1 vssd1 vccd1 vccd1 _18583_/A sky130_fd_sc_hd__and3_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _17533_/A vssd1 vssd1 vccd1 vccd1 _25843_/D sky130_fd_sc_hd__clkbuf_1
X_14745_ _14743_/X _26543_/Q _14757_/S vssd1 vssd1 vccd1 vccd1 _14746_/A sky130_fd_sc_hd__mux2_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17464_ _17463_/X _25823_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17465_/A sky130_fd_sc_hd__mux2_1
X_14676_ _26567_/Q _14671_/X _14666_/X _14675_/Y vssd1 vssd1 vccd1 vccd1 _26567_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19203_ _19338_/A vssd1 vssd1 vccd1 vccd1 _19203_/X sky130_fd_sc_hd__buf_2
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16415_ _16734_/B vssd1 vssd1 vccd1 vccd1 _16708_/A sky130_fd_sc_hd__clkbuf_2
X_13627_ _13897_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13627_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17395_ input74/X vssd1 vssd1 vccd1 vccd1 _20796_/A sky130_fd_sc_hd__inv_2
XFILLER_9_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19134_ _19132_/X _19133_/X _19499_/S vssd1 vssd1 vccd1 vccd1 _19134_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16346_ _16862_/B _16347_/B vssd1 vssd1 vccd1 vccd1 _16864_/B sky130_fd_sc_hd__xor2_1
XFILLER_160_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater85 _27296_/CLK vssd1 vssd1 vccd1 vccd1 _27423_/CLK sky130_fd_sc_hd__clkbuf_1
X_13558_ _13558_/A vssd1 vssd1 vccd1 vccd1 _13558_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater96 _26030_/CLK vssd1 vssd1 vccd1 vccd1 _25935_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19065_ _26691_/Q _26659_/Q _26627_/Q _26595_/Q _18908_/X _18909_/X vssd1 vssd1 vccd1
+ vccd1 _19066_/B sky130_fd_sc_hd__mux4_2
XFILLER_157_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16277_ _16277_/A _16277_/B vssd1 vssd1 vccd1 vccd1 _16277_/Y sky130_fd_sc_hd__nor2_1
X_13489_ _16536_/A vssd1 vssd1 vccd1 vccd1 _13889_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18016_ _27597_/Q vssd1 vssd1 vccd1 vccd1 _18016_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15228_ _14763_/X _26345_/Q _15234_/S vssd1 vssd1 vccd1 vccd1 _15229_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15159_ _15159_/A vssd1 vssd1 vccd1 vccd1 _26376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19967_ _19967_/A vssd1 vssd1 vccd1 vccd1 _19967_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18918_ _24403_/A _18916_/X _24405_/A vssd1 vssd1 vccd1 vccd1 _18918_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19898_ _19898_/A vssd1 vssd1 vccd1 vccd1 _19898_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18849_ _18775_/X _18848_/X _18785_/X vssd1 vssd1 vccd1 vccd1 _18849_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21860_ _21860_/A vssd1 vssd1 vccd1 vccd1 _21860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20811_ _20811_/A vssd1 vssd1 vccd1 vccd1 _20811_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21791_ _21777_/X _21778_/X _21779_/X _21780_/X _21781_/X _21782_/X vssd1 vssd1 vccd1
+ vccd1 _21792_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23530_ _24844_/A _27200_/Q _23542_/S vssd1 vssd1 vccd1 vccd1 _23531_/B sky130_fd_sc_hd__mux2_1
XFILLER_196_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20742_ _20758_/A vssd1 vssd1 vccd1 vccd1 _20742_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23461_ _25132_/A vssd1 vssd1 vccd1 vccd1 _23461_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20673_ _20673_/A vssd1 vssd1 vccd1 vccd1 _20673_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25200_ _27700_/Q _25184_/X _25199_/Y _25175_/X vssd1 vssd1 vccd1 vccd1 _27700_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22412_ _22412_/A vssd1 vssd1 vccd1 vccd1 _22412_/X sky130_fd_sc_hd__clkbuf_1
X_26180_ _19947_/X _26180_/D vssd1 vssd1 vccd1 vccd1 _26180_/Q sky130_fd_sc_hd__dfxtp_1
X_23392_ _24754_/A _27241_/Q _27244_/Q _24763_/A _23391_/X vssd1 vssd1 vccd1 vccd1
+ _23393_/D sky130_fd_sc_hd__a221o_1
XFILLER_192_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25131_ _25139_/A _25131_/B vssd1 vssd1 vccd1 vccd1 _25131_/Y sky130_fd_sc_hd__nand2_1
X_22343_ _22331_/X _22332_/X _22333_/X _22334_/X _22335_/X _22336_/X vssd1 vssd1 vccd1
+ vccd1 _22344_/A sky130_fd_sc_hd__mux4_1
XFILLER_137_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25062_ _27836_/Q _27140_/Q _25885_/Q _25853_/Q _25061_/X _25035_/X vssd1 vssd1 vccd1
+ vccd1 _25062_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_806 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22274_ _22274_/A vssd1 vssd1 vccd1 vccd1 _22274_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24013_ _23990_/X _24011_/X _24012_/X _24005_/X vssd1 vssd1 vccd1 vccd1 _27297_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21225_ _21211_/X _21212_/X _21213_/X _21214_/X _21216_/X _21218_/X vssd1 vssd1 vccd1
+ vccd1 _21226_/A sky130_fd_sc_hd__mux4_1
XFILLER_176_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21156_ _21156_/A vssd1 vssd1 vccd1 vccd1 _21156_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20107_ _20107_/A vssd1 vssd1 vccd1 vccd1 _20107_/X sky130_fd_sc_hd__clkbuf_1
X_25964_ _27326_/CLK _25964_/D vssd1 vssd1 vccd1 vccd1 _25964_/Q sky130_fd_sc_hd__dfxtp_1
X_21087_ _21077_/X _21078_/X _21079_/X _21080_/X _21081_/X _21082_/X vssd1 vssd1 vccd1
+ vccd1 _21088_/A sky130_fd_sc_hd__mux4_1
XFILLER_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27703_ _27703_/CLK _27703_/D vssd1 vssd1 vccd1 vccd1 _27703_/Q sky130_fd_sc_hd__dfxtp_1
X_24915_ _27659_/Q _24909_/X _24913_/Y _24914_/X vssd1 vssd1 vccd1 vccd1 _27659_/D
+ sky130_fd_sc_hd__o211a_1
X_20038_ _20028_/X _20029_/X _20030_/X _20031_/X _20032_/X _20033_/X vssd1 vssd1 vccd1
+ vccd1 _20039_/A sky130_fd_sc_hd__mux4_1
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25895_ _25895_/CLK _25895_/D vssd1 vssd1 vccd1 vccd1 _25895_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27634_ _27636_/CLK _27634_/D vssd1 vssd1 vccd1 vccd1 _27634_/Q sky130_fd_sc_hd__dfxtp_1
X_24846_ _24863_/A _24846_/B vssd1 vssd1 vccd1 vccd1 _24846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27565_ _27569_/CLK _27565_/D vssd1 vssd1 vccd1 vccd1 _27565_/Q sky130_fd_sc_hd__dfxtp_1
X_24777_ _27624_/Q _24771_/X _24776_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _27624_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ _21981_/X _21982_/X _21983_/X _21984_/X _21985_/X _21986_/X vssd1 vssd1 vccd1
+ vccd1 _21990_/A sky130_fd_sc_hd__mux4_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14530_/A vssd1 vssd1 vccd1 vccd1 _14530_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26516_ _21118_/X _26516_/D vssd1 vssd1 vccd1 vccd1 _26516_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23728_ _23728_/A vssd1 vssd1 vccd1 vccd1 _27266_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27496_ _27527_/CLK _27496_/D vssd1 vssd1 vccd1 vccd1 _27496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14461_ _16536_/A vssd1 vssd1 vccd1 vccd1 _15730_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26447_ _20880_/X _26447_/D vssd1 vssd1 vccd1 vccd1 _26447_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23659_ _24835_/B _27236_/Q _23661_/S vssd1 vssd1 vccd1 vccd1 _23660_/A sky130_fd_sc_hd__mux2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16200_ _16345_/A _16200_/B _16756_/A _16326_/A vssd1 vssd1 vccd1 vccd1 _16358_/A
+ sky130_fd_sc_hd__or4_1
X_13412_ _26973_/Q _13411_/X _13415_/S vssd1 vssd1 vccd1 vccd1 _13413_/A sky130_fd_sc_hd__mux2_1
X_17180_ _17155_/X _17180_/B vssd1 vssd1 vccd1 vccd1 _17180_/X sky130_fd_sc_hd__and2b_1
X_14392_ _14441_/A vssd1 vssd1 vccd1 vccd1 _14392_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26378_ _20633_/X _26378_/D vssd1 vssd1 vccd1 vccd1 _26378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _16264_/B _16296_/B _26070_/Q vssd1 vssd1 vccd1 vccd1 _16131_/X sky130_fd_sc_hd__or3b_1
X_25329_ _25329_/A _25329_/B _25329_/C _25329_/D vssd1 vssd1 vccd1 vccd1 _25329_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_6_611 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ _13343_/A vssd1 vssd1 vccd1 vccd1 _26995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16062_ _16062_/A _16062_/B vssd1 vssd1 vccd1 vccd1 _16063_/D sky130_fd_sc_hd__or2_1
XFILLER_170_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _27022_/Q _13122_/X _13280_/S vssd1 vssd1 vccd1 vccd1 _13275_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15013_ _15751_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _15013_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19821_ _19821_/A vssd1 vssd1 vccd1 vccd1 _19821_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19752_ _19800_/A vssd1 vssd1 vccd1 vccd1 _19752_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16964_ _24633_/A _24522_/A _16982_/C _16963_/X vssd1 vssd1 vccd1 vccd1 _16967_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18703_ _18703_/A vssd1 vssd1 vccd1 vccd1 _26014_/D sky130_fd_sc_hd__clkbuf_1
X_15915_ _15918_/A vssd1 vssd1 vccd1 vccd1 _15915_/Y sky130_fd_sc_hd__inv_2
X_19683_ _19715_/A vssd1 vssd1 vccd1 vccd1 _19683_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16895_ _24262_/A _24249_/A _24256_/A _24232_/A vssd1 vssd1 vccd1 vccd1 _16895_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _18634_/A vssd1 vssd1 vccd1 vccd1 _25983_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _15846_/A vssd1 vssd1 vccd1 vccd1 _26078_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18565_ _18565_/A vssd1 vssd1 vccd1 vccd1 _25974_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _15777_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15777_/Y sky130_fd_sc_hd__nor2_1
X_12989_ _13000_/A vssd1 vssd1 vccd1 vccd1 _12998_/B sky130_fd_sc_hd__clkbuf_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17516_ _17516_/A vssd1 vssd1 vccd1 vccd1 _25839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14728_ _14811_/S vssd1 vssd1 vccd1 vccd1 _14741_/S sky130_fd_sc_hd__clkbuf_2
X_18496_ _26837_/Q _26805_/Q _26773_/Q _26741_/Q _17832_/X _18380_/X vssd1 vssd1 vccd1
+ vccd1 _18496_/X sky130_fd_sc_hd__mux4_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14659_ _15732_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17447_ _27415_/Q vssd1 vssd1 vccd1 vccd1 _17447_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17378_ _17378_/A vssd1 vssd1 vccd1 vccd1 _27946_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_158_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19117_ _26949_/Q _26917_/Q _26885_/Q _26853_/Q _19044_/X _19116_/X vssd1 vssd1 vccd1
+ vccd1 _19117_/X sky130_fd_sc_hd__mux4_2
XFILLER_145_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16329_ _16862_/A _16200_/B _16369_/A vssd1 vssd1 vccd1 vccd1 _16336_/B sky130_fd_sc_hd__o21a_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _19041_/X _19043_/X _19047_/X _19022_/X _19023_/X vssd1 vssd1 vccd1 vccd1
+ _19059_/B sky130_fd_sc_hd__a221o_1
XFILLER_145_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21010_ _21042_/A vssd1 vssd1 vccd1 vccd1 _21010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_415 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22961_ _22961_/A vssd1 vssd1 vccd1 vccd1 _23030_/A sky130_fd_sc_hd__clkbuf_4
X_24700_ _24700_/A vssd1 vssd1 vccd1 vccd1 _24700_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21912_ _21912_/A vssd1 vssd1 vccd1 vccd1 _21912_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25680_ _25680_/A vssd1 vssd1 vccd1 vccd1 _25680_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22892_ _22957_/A vssd1 vssd1 vccd1 vccd1 _22892_/X sky130_fd_sc_hd__clkbuf_1
X_24631_ _24631_/A _24631_/B vssd1 vssd1 vccd1 vccd1 _24632_/A sky130_fd_sc_hd__and2_1
XFILLER_83_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21843_ _22015_/A vssd1 vssd1 vccd1 vccd1 _21911_/A sky130_fd_sc_hd__buf_2
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27350_ _27350_/CLK _27350_/D vssd1 vssd1 vccd1 vccd1 _27350_/Q sky130_fd_sc_hd__dfxtp_2
X_24562_ _24562_/A vssd1 vssd1 vccd1 vccd1 _27542_/D sky130_fd_sc_hd__clkbuf_1
X_21774_ _21774_/A vssd1 vssd1 vccd1 vccd1 _21774_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26301_ _20369_/X _26301_/D vssd1 vssd1 vccd1 vccd1 _26301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23513_ _25977_/Q _27196_/Q _23525_/S vssd1 vssd1 vccd1 vccd1 _23514_/B sky130_fd_sc_hd__mux2_1
X_27281_ _27418_/CLK _27281_/D vssd1 vssd1 vccd1 vccd1 _27281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20725_ _20773_/A vssd1 vssd1 vccd1 vccd1 _20725_/X sky130_fd_sc_hd__clkbuf_1
X_24493_ _27584_/Q _24493_/B vssd1 vssd1 vccd1 vccd1 _24629_/B sky130_fd_sc_hd__nor2_1
X_26232_ _20125_/X _26232_/D vssd1 vssd1 vccd1 vccd1 _26232_/Q sky130_fd_sc_hd__dfxtp_1
X_23444_ input40/X _23442_/X _23443_/X _23434_/X vssd1 vssd1 vccd1 vccd1 _27171_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20656_ _20672_/A vssd1 vssd1 vccd1 vccd1 _20656_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26163_ _19879_/X _26163_/D vssd1 vssd1 vccd1 vccd1 _26163_/Q sky130_fd_sc_hd__dfxtp_1
X_23375_ _27757_/Q _23334_/Y _27261_/Q _24808_/A _23374_/X vssd1 vssd1 vccd1 vccd1
+ _23410_/B sky130_fd_sc_hd__a221o_1
X_20587_ _20587_/A vssd1 vssd1 vccd1 vccd1 _20587_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25114_ _27689_/Q _25112_/X _25113_/Y _23498_/X vssd1 vssd1 vccd1 vccd1 _27689_/D
+ sky130_fd_sc_hd__o211a_1
X_22326_ _22326_/A vssd1 vssd1 vccd1 vccd1 _22326_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26094_ _19636_/X _26094_/D vssd1 vssd1 vccd1 vccd1 _26094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25045_ _25920_/Q _25986_/Q _25819_/Q _26018_/Q _25009_/X _25027_/X vssd1 vssd1 vccd1
+ vccd1 _25045_/X sky130_fd_sc_hd__mux4_1
X_22257_ _22245_/X _22246_/X _22247_/X _22248_/X _22249_/X _22250_/X vssd1 vssd1 vccd1
+ vccd1 _22258_/A sky130_fd_sc_hd__mux4_1
XFILLER_152_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21208_ _21208_/A vssd1 vssd1 vccd1 vccd1 _21208_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22188_ _22188_/A vssd1 vssd1 vccd1 vccd1 _22188_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_437 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21139_ _21125_/X _21126_/X _21127_/X _21128_/X _21130_/X _21132_/X vssd1 vssd1 vccd1
+ vccd1 _21140_/A sky130_fd_sc_hd__mux4_1
XFILLER_63_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26996_ _22794_/X _26996_/D vssd1 vssd1 vccd1 vccd1 _26996_/Q sky130_fd_sc_hd__dfxtp_1
X_13961_ _14433_/A vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__buf_2
XFILLER_120_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25947_ _27312_/CLK _25947_/D vssd1 vssd1 vccd1 vccd1 _25947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15700_ _26137_/Q _15040_/X _15697_/X _15699_/Y vssd1 vssd1 vccd1 vccd1 _26137_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16680_ _16751_/B vssd1 vssd1 vccd1 vccd1 _16681_/B sky130_fd_sc_hd__inv_2
X_13892_ _26829_/Q _13880_/X _13886_/X _13891_/Y vssd1 vssd1 vccd1 vccd1 _26829_/D
+ sky130_fd_sc_hd__a31o_1
X_25878_ _25878_/CLK _25878_/D vssd1 vssd1 vccd1 vccd1 _25878_/Q sky130_fd_sc_hd__dfxtp_1
X_27617_ _27617_/CLK _27617_/D vssd1 vssd1 vccd1 vccd1 _27617_/Q sky130_fd_sc_hd__dfxtp_1
X_24829_ _24829_/A vssd1 vssd1 vccd1 vccd1 _27642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _15631_/A vssd1 vssd1 vccd1 vccd1 _26167_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _18348_/X _18349_/X _18395_/A vssd1 vssd1 vccd1 vccd1 _18350_/X sky130_fd_sc_hd__mux2_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _26197_/Q _14724_/A _15562_/S vssd1 vssd1 vccd1 vccd1 _15563_/A sky130_fd_sc_hd__mux2_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27548_ _27668_/CLK _27548_/D vssd1 vssd1 vccd1 vccd1 _27548_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _25936_/Q _26002_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17302_/B sky130_fd_sc_hd__mux2_1
X_14513_ _26624_/Q _14496_/X _14510_/X _14512_/Y vssd1 vssd1 vccd1 vccd1 _26624_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18281_ _18279_/X _18280_/X _18211_/X vssd1 vssd1 vccd1 vccd1 _18281_/X sky130_fd_sc_hd__o21a_1
X_27479_ _27572_/CLK _27479_/D vssd1 vssd1 vccd1 vccd1 _27479_/Q sky130_fd_sc_hd__dfxtp_1
X_15493_ _13086_/X _26228_/Q _15501_/S vssd1 vssd1 vccd1 vccd1 _15494_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17232_ _17181_/X _17231_/X _17220_/X vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__a21bo_1
X_14444_ _26643_/Q _14441_/X _14437_/X _14443_/Y vssd1 vssd1 vccd1 vccd1 _26643_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17163_ _17161_/X _17162_/X _17174_/S vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__mux2_2
XFILLER_122_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ _26665_/Q _14365_/X _14371_/X _14374_/Y vssd1 vssd1 vccd1 vccd1 _26665_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _16191_/B vssd1 vssd1 vccd1 vccd1 _16235_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_155_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _27000_/Q _13325_/X _13335_/S vssd1 vssd1 vccd1 vccd1 _13327_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17094_ _17303_/A vssd1 vssd1 vccd1 vccd1 _17094_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16045_ _27477_/Q _27373_/Q vssd1 vssd1 vccd1 vccd1 _16045_/X sky130_fd_sc_hd__xor2_1
X_13257_ _13257_/A vssd1 vssd1 vccd1 vccd1 _27030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13188_ _27343_/Q _13017_/A _13025_/A _27311_/Q _13187_/X vssd1 vssd1 vccd1 vccd1
+ _16230_/A sky130_fd_sc_hd__a221o_1
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19804_ _19796_/X _19797_/X _19798_/X _19799_/X _19800_/X _19801_/X vssd1 vssd1 vccd1
+ vccd1 _19805_/A sky130_fd_sc_hd__mux4_1
XFILLER_150_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17996_ _18462_/A vssd1 vssd1 vccd1 vccd1 _17996_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19735_ _19735_/A vssd1 vssd1 vccd1 vccd1 _19735_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16947_ _27577_/Q _16947_/B vssd1 vssd1 vccd1 vccd1 _24640_/A sky130_fd_sc_hd__and2_1
XFILLER_38_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19666_ _19714_/A vssd1 vssd1 vccd1 vccd1 _19666_/X sky130_fd_sc_hd__clkbuf_2
X_16878_ _16599_/Y _16878_/B vssd1 vssd1 vccd1 vccd1 _16879_/C sky130_fd_sc_hd__and2b_1
XFILLER_65_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18617_ _24828_/A _18606_/X _24825_/A vssd1 vssd1 vccd1 vccd1 _18617_/Y sky130_fd_sc_hd__o21ai_1
X_15829_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15838_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19597_ _19589_/X _19590_/X _19591_/X _19592_/X _19593_/X _19594_/X vssd1 vssd1 vccd1
+ vccd1 _19598_/A sky130_fd_sc_hd__mux4_1
XFILLER_92_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18548_ _27823_/Q _26584_/Q _26456_/Q _26136_/Q _17789_/X _18425_/X vssd1 vssd1 vccd1
+ vccd1 _18548_/X sky130_fd_sc_hd__mux4_1
X_18479_ _18479_/A vssd1 vssd1 vccd1 vccd1 _18479_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20510_ _20496_/X _20497_/X _20498_/X _20499_/X _20500_/X _20501_/X vssd1 vssd1 vccd1
+ vccd1 _20511_/A sky130_fd_sc_hd__mux4_1
X_21490_ _21490_/A vssd1 vssd1 vccd1 vccd1 _21490_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20441_ _20441_/A vssd1 vssd1 vccd1 vccd1 _20441_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23160_ _23160_/A vssd1 vssd1 vccd1 vccd1 _27119_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20372_ _20354_/X _20357_/X _20360_/X _20363_/X _20364_/X _20365_/X vssd1 vssd1 vccd1
+ vccd1 _20373_/A sky130_fd_sc_hd__mux4_1
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22111_ _22457_/A vssd1 vssd1 vccd1 vccd1 _22176_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23091_ _23091_/A vssd1 vssd1 vccd1 vccd1 _27089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22042_ _22042_/A vssd1 vssd1 vccd1 vccd1 _22042_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26850_ _22290_/X _26850_/D vssd1 vssd1 vccd1 vccd1 _26850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25801_ _17517_/X _27855_/Q _25801_/S vssd1 vssd1 vccd1 vccd1 _25802_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26781_ _22044_/X _26781_/D vssd1 vssd1 vccd1 vccd1 _26781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23993_ _27785_/Q vssd1 vssd1 vccd1 vccd1 _23993_/X sky130_fd_sc_hd__buf_2
X_25732_ _25732_/A vssd1 vssd1 vccd1 vccd1 _25732_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22944_ _22944_/A vssd1 vssd1 vccd1 vccd1 _22944_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25663_ _25654_/X _25656_/X _25658_/X _25660_/X _25661_/X _25662_/X vssd1 vssd1 vccd1
+ vccd1 _25664_/A sky130_fd_sc_hd__mux4_1
X_22875_ _22961_/A vssd1 vssd1 vccd1 vccd1 _22944_/A sky130_fd_sc_hd__buf_2
XFILLER_37_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27402_ _27402_/CLK _27402_/D vssd1 vssd1 vccd1 vccd1 _27402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24614_ _27666_/Q _24620_/B vssd1 vssd1 vccd1 vccd1 _24615_/A sky130_fd_sc_hd__and2_1
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21826_ _21826_/A vssd1 vssd1 vccd1 vccd1 _21826_/X sky130_fd_sc_hd__clkbuf_1
X_25594_ _25572_/X _25582_/X _25583_/X _24952_/B _25584_/X vssd1 vssd1 vccd1 vccd1
+ _25594_/X sky130_fd_sc_hd__o311a_1
XFILLER_93_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27333_ _27333_/CLK _27333_/D vssd1 vssd1 vccd1 vccd1 _27333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24545_ _24534_/X _24392_/A _24545_/S vssd1 vssd1 vccd1 vccd1 _24546_/B sky130_fd_sc_hd__mux2_1
X_21757_ _22015_/A vssd1 vssd1 vccd1 vccd1 _21825_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20708_ _20708_/A vssd1 vssd1 vccd1 vccd1 _20773_/A sky130_fd_sc_hd__buf_2
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27264_ _27264_/CLK _27264_/D vssd1 vssd1 vccd1 vccd1 _27264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24476_ _27635_/Q _24478_/B vssd1 vssd1 vccd1 vccd1 _24477_/A sky130_fd_sc_hd__and2_1
X_21688_ _21688_/A vssd1 vssd1 vccd1 vccd1 _21688_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26215_ _20067_/X _26215_/D vssd1 vssd1 vccd1 vccd1 _26215_/Q sky130_fd_sc_hd__dfxtp_1
X_23427_ _27165_/Q _23430_/B vssd1 vssd1 vccd1 vccd1 _23427_/X sky130_fd_sc_hd__or2_1
X_20639_ _20687_/A vssd1 vssd1 vccd1 vccd1 _20639_/X sky130_fd_sc_hd__clkbuf_1
X_27195_ _27196_/CLK _27195_/D vssd1 vssd1 vccd1 vccd1 _27195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ _14166_/A vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26146_ _19823_/X _26146_/D vssd1 vssd1 vccd1 vccd1 _26146_/Q sky130_fd_sc_hd__dfxtp_1
X_23358_ _24759_/A _27243_/Q _27260_/Q _24806_/A vssd1 vssd1 vccd1 vccd1 _23358_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _14740_/A vssd1 vssd1 vccd1 vccd1 _13111_/X sky130_fd_sc_hd__buf_2
X_22309_ _22299_/X _22300_/X _22301_/X _22302_/X _22303_/X _22304_/X vssd1 vssd1 vccd1
+ vccd1 _22310_/A sky130_fd_sc_hd__mux4_1
XFILLER_166_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14091_ _14356_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14091_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26077_ _19584_/X _26077_/D vssd1 vssd1 vccd1 vccd1 _26077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23289_ _23280_/Y input41/X _27726_/Q _23288_/Y vssd1 vssd1 vccd1 vccd1 _23293_/C
+ sky130_fd_sc_hd__o22ai_1
XFILLER_152_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13042_ _16014_/B vssd1 vssd1 vccd1 vccd1 _15045_/B sky130_fd_sc_hd__clkbuf_2
X_25028_ _25918_/Q _25984_/Q _25817_/Q _26016_/Q _25009_/X _25027_/X vssd1 vssd1 vccd1
+ vccd1 _25028_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17850_ _17924_/A vssd1 vssd1 vccd1 vccd1 _18405_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_61_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16801_ _16801_/A _16822_/A vssd1 vssd1 vccd1 vccd1 _16801_/X sky130_fd_sc_hd__or2_1
XFILLER_120_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17781_ _18360_/A vssd1 vssd1 vccd1 vccd1 _18458_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_120_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14993_ _26446_/Q _14988_/X _14989_/X _14992_/Y vssd1 vssd1 vccd1 vccd1 _26446_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26979_ _22734_/X _26979_/D vssd1 vssd1 vccd1 vccd1 _26979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19520_ _27822_/Q _26583_/Q _26455_/Q _26135_/Q _19414_/X _18831_/X vssd1 vssd1 vccd1
+ vccd1 _19520_/X sky130_fd_sc_hd__mux4_1
X_16732_ _16732_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16732_/Y sky130_fd_sc_hd__xnor2_1
X_13944_ _14060_/B vssd1 vssd1 vccd1 vccd1 _13944_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19451_ _19451_/A vssd1 vssd1 vccd1 vccd1 _26067_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13875_ _26836_/Q _13865_/X _13873_/X _13874_/Y vssd1 vssd1 vccd1 vccd1 _26836_/D
+ sky130_fd_sc_hd__a31o_1
X_16663_ _16626_/X _16658_/Y _16659_/Y _16662_/X _16619_/X vssd1 vssd1 vccd1 vccd1
+ _24253_/A sky130_fd_sc_hd__a32o_1
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18402_ _27816_/Q _26577_/Q _26449_/Q _26129_/Q _18401_/X _18267_/X vssd1 vssd1 vccd1
+ vccd1 _18402_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15614_ _15614_/A vssd1 vssd1 vccd1 vccd1 _26174_/D sky130_fd_sc_hd__clkbuf_1
X_19382_ _19382_/A vssd1 vssd1 vccd1 vccd1 _26064_/D sky130_fd_sc_hd__clkbuf_1
X_16594_ _16594_/A vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18333_ _18398_/A _18333_/B _18333_/C vssd1 vssd1 vccd1 vccd1 _18334_/A sky130_fd_sc_hd__and3_1
XFILLER_72_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15545_ _13228_/X _26204_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15546_/A sky130_fd_sc_hd__mux2_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15476_ _15476_/A vssd1 vssd1 vccd1 vccd1 _26235_/D sky130_fd_sc_hd__clkbuf_1
X_18264_ _18264_/A _18264_/B _18264_/C vssd1 vssd1 vccd1 vccd1 _18265_/A sky130_fd_sc_hd__and3_1
X_17215_ _27843_/Q _27147_/Q _25892_/Q _25860_/Q _17203_/X _17191_/X vssd1 vssd1 vccd1
+ vccd1 _17215_/X sky130_fd_sc_hd__mux4_1
X_14427_ _26647_/Q _14421_/X _14416_/X _14426_/Y vssd1 vssd1 vccd1 vccd1 _26647_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18195_ _27807_/Q _26568_/Q _26440_/Q _26120_/Q _18099_/X _18126_/X vssd1 vssd1 vccd1
+ vccd1 _18195_/X sky130_fd_sc_hd__mux4_2
X_14358_ _14398_/A vssd1 vssd1 vccd1 vccd1 _14358_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17146_ _17094_/X _17146_/B vssd1 vssd1 vccd1 vccd1 _17146_/X sky130_fd_sc_hd__and2b_1
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13309_ _27006_/Q _13216_/X _13313_/S vssd1 vssd1 vccd1 vccd1 _13310_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17077_ _17075_/X _17076_/X _17113_/S vssd1 vssd1 vccd1 vccd1 _17077_/X sky130_fd_sc_hd__mux2_1
X_14289_ _14376_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16028_ _16287_/A vssd1 vssd1 vccd1 vccd1 _16144_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17979_ _17979_/A _17978_/X vssd1 vssd1 vccd1 vccd1 _17979_/X sky130_fd_sc_hd__or2b_1
XFILLER_85_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19718_ _19710_/X _19711_/X _19712_/X _19713_/X _19714_/X _19715_/X vssd1 vssd1 vccd1
+ vccd1 _19719_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20990_ _20990_/A vssd1 vssd1 vccd1 vccd1 _20990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19649_ _19649_/A vssd1 vssd1 vccd1 vccd1 _19649_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22660_ _22660_/A vssd1 vssd1 vccd1 vccd1 _22660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21611_ _21599_/X _21600_/X _21601_/X _21602_/X _21603_/X _21604_/X vssd1 vssd1 vccd1
+ vccd1 _21612_/A sky130_fd_sc_hd__mux4_1
X_22591_ _22577_/X _22578_/X _22579_/X _22580_/X _22581_/X _22582_/X vssd1 vssd1 vccd1
+ vccd1 _22592_/A sky130_fd_sc_hd__mux4_1
XFILLER_139_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24330_ _24330_/A vssd1 vssd1 vccd1 vccd1 _24339_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_194_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21542_ _21542_/A vssd1 vssd1 vccd1 vccd1 _21542_/X sky130_fd_sc_hd__clkbuf_1
X_24261_ _24261_/A _24264_/B vssd1 vssd1 vccd1 vccd1 _27403_/D sky130_fd_sc_hd__nor2_1
XFILLER_193_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21473_ _21459_/X _21460_/X _21461_/X _21462_/X _21463_/X _21464_/X vssd1 vssd1 vccd1
+ vccd1 _21474_/A sky130_fd_sc_hd__mux4_1
XFILLER_14_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26000_ _26001_/CLK _26000_/D vssd1 vssd1 vccd1 vccd1 _26000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23212_ _23212_/A vssd1 vssd1 vccd1 vccd1 _27142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20424_ _20424_/A vssd1 vssd1 vccd1 vccd1 _20424_/X sky130_fd_sc_hd__clkbuf_1
X_24192_ _24192_/A vssd1 vssd1 vccd1 vccd1 _27366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23143_ _27112_/Q _17721_/X _23143_/S vssd1 vssd1 vccd1 vccd1 _23144_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20355_ _25655_/A vssd1 vssd1 vccd1 vccd1 _20704_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27951_ _27951_/A _15924_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
X_23074_ _23074_/A vssd1 vssd1 vccd1 vccd1 _27081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20286_ _20334_/A vssd1 vssd1 vccd1 vccd1 _20286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22025_ _22016_/X _22018_/X _22020_/X _22022_/X _22023_/X _22024_/X vssd1 vssd1 vccd1
+ vccd1 _22026_/A sky130_fd_sc_hd__mux4_1
X_26902_ _22466_/X _26902_/D vssd1 vssd1 vccd1 vccd1 _26902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26833_ _22226_/X _26833_/D vssd1 vssd1 vccd1 vccd1 _26833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26764_ _21980_/X _26764_/D vssd1 vssd1 vccd1 vccd1 _26764_/Q sky130_fd_sc_hd__dfxtp_1
X_23976_ _27786_/Q vssd1 vssd1 vccd1 vccd1 _23976_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22927_ _22943_/A vssd1 vssd1 vccd1 vccd1 _22927_/X sky130_fd_sc_hd__clkbuf_2
X_25715_ _25705_/X _25706_/X _25707_/X _25708_/X _25709_/X _25710_/X vssd1 vssd1 vccd1
+ vccd1 _25716_/A sky130_fd_sc_hd__mux4_1
X_26695_ _21748_/X _26695_/D vssd1 vssd1 vccd1 vccd1 _26695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ _26911_/Q _13653_/X _13656_/X _13659_/Y vssd1 vssd1 vccd1 vccd1 _26911_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22858_ _22858_/A vssd1 vssd1 vccd1 vccd1 _22858_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25646_ _25646_/A vssd1 vssd1 vccd1 vccd1 _25646_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21809_ _21825_/A vssd1 vssd1 vccd1 vccd1 _21809_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13859_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13591_/Y sky130_fd_sc_hd__nor2_1
X_25577_ _24267_/A _25440_/X _25442_/X _24937_/B _24384_/A vssd1 vssd1 vccd1 vccd1
+ _25577_/X sky130_fd_sc_hd__o311a_1
XFILLER_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22789_ _22961_/A vssd1 vssd1 vccd1 vccd1 _22858_/A sky130_fd_sc_hd__clkbuf_2
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _26299_/Q _13417_/X _15332_/S vssd1 vssd1 vccd1 vccd1 _15331_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24528_ _24631_/A _24528_/B vssd1 vssd1 vccd1 vccd1 _24529_/A sky130_fd_sc_hd__and2_1
X_27316_ _27331_/CLK _27316_/D vssd1 vssd1 vccd1 vccd1 _27316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _15261_/A vssd1 vssd1 vccd1 vccd1 _26330_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24459_ _27627_/Q _24467_/B vssd1 vssd1 vccd1 vccd1 _24460_/A sky130_fd_sc_hd__and2_1
X_27247_ _27263_/CLK _27247_/D vssd1 vssd1 vccd1 vccd1 _27247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ _14225_/A vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17000_ _25811_/Q _26010_/Q _17061_/A vssd1 vssd1 vccd1 vccd1 _17000_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1165 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27178_ _27180_/CLK _27178_/D vssd1 vssd1 vccd1 vccd1 _27178_/Q sky130_fd_sc_hd__dfxtp_1
X_15192_ _15260_/S vssd1 vssd1 vccd1 vccd1 _15201_/S sky130_fd_sc_hd__buf_2
XFILLER_126_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_412 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _25824_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14408_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _14143_/Y sky130_fd_sc_hd__nor2_1
X_26129_ _19763_/X _26129_/D vssd1 vssd1 vccd1 vccd1 _26129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14074_ _14340_/A _14085_/B vssd1 vssd1 vccd1 vccd1 _14074_/Y sky130_fd_sc_hd__nor2_1
X_18951_ _26142_/Q _26078_/Q _27006_/Q _26974_/Q _18882_/X _18950_/X vssd1 vssd1 vccd1
+ vccd1 _18952_/B sky130_fd_sc_hd__mux4_1
XFILLER_180_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17902_ _26524_/Q _26492_/Q _26460_/Q _27036_/Q _17899_/X _17901_/X vssd1 vssd1 vccd1
+ vccd1 _17902_/X sky130_fd_sc_hd__mux4_1
X_13025_ _13025_/A vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18882_ _19165_/A vssd1 vssd1 vccd1 vccd1 _18882_/X sky130_fd_sc_hd__buf_2
XFILLER_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17833_ _17900_/A vssd1 vssd1 vccd1 vccd1 _18408_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17764_ _25939_/Q _17763_/X _17770_/S vssd1 vssd1 vccd1 vccd1 _17765_/A sky130_fd_sc_hd__mux2_1
X_14976_ _15029_/A vssd1 vssd1 vccd1 vccd1 _14976_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19503_ _18929_/X _19502_/X _18932_/X vssd1 vssd1 vccd1 vccd1 _19503_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16715_ _16852_/A _16715_/B _16715_/C _16737_/B vssd1 vssd1 vccd1 vccd1 _16731_/A
+ sky130_fd_sc_hd__or4_1
X_13927_ _26816_/Q _13919_/X _13925_/X _13926_/Y vssd1 vssd1 vccd1 vccd1 _26816_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_484 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17695_ _17695_/A vssd1 vssd1 vccd1 vccd1 _25917_/D sky130_fd_sc_hd__clkbuf_1
X_19434_ _26963_/Q _26931_/Q _26899_/Q _26867_/Q _19343_/X _19412_/X vssd1 vssd1 vccd1
+ vccd1 _19434_/X sky130_fd_sc_hd__mux4_1
X_16646_ _25909_/Q _16646_/B vssd1 vssd1 vccd1 vccd1 _16647_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _26841_/Q _13844_/X _13855_/X _13857_/Y vssd1 vssd1 vccd1 vccd1 _26841_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19365_ _26960_/Q _26928_/Q _26896_/Q _26864_/Q _19061_/X _18920_/X vssd1 vssd1 vccd1
+ vccd1 _19365_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16577_ _16833_/A _16577_/B vssd1 vssd1 vccd1 vccd1 _16585_/B sky130_fd_sc_hd__xnor2_1
X_13789_ _26865_/Q _13778_/X _13780_/X _13788_/Y vssd1 vssd1 vccd1 vccd1 _26865_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18316_ _26701_/Q _26669_/Q _26637_/Q _26605_/Q _18177_/X _18249_/X vssd1 vssd1 vccd1
+ vccd1 _18318_/A sky130_fd_sc_hd__mux4_2
X_15528_ _13179_/X _26212_/Q _15534_/S vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__mux2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19296_ _19294_/X _19295_/X _19296_/S vssd1 vssd1 vccd1 vccd1 _19296_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ _18243_/X _18245_/X _18378_/S vssd1 vssd1 vccd1 vccd1 _18247_/X sky130_fd_sc_hd__mux2_1
X_15459_ _15459_/A vssd1 vssd1 vccd1 vccd1 _26243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18178_ _26695_/Q _26663_/Q _26631_/Q _26599_/Q _18177_/X _18106_/X vssd1 vssd1 vccd1
+ vccd1 _18179_/A sky130_fd_sc_hd__mux4_1
XFILLER_128_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_591 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17129_ _17129_/A vssd1 vssd1 vccd1 vccd1 _27925_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_171_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20140_ _20130_/X _20131_/X _20132_/X _20133_/X _20134_/X _20135_/X vssd1 vssd1 vccd1
+ vccd1 _20141_/A sky130_fd_sc_hd__mux4_1
XFILLER_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ _20071_/A vssd1 vssd1 vccd1 vccd1 _20071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater320 _27511_/CLK vssd1 vssd1 vccd1 vccd1 _27515_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater331 _27774_/CLK vssd1 vssd1 vccd1 vccd1 _27716_/CLK sky130_fd_sc_hd__clkbuf_1
X_23830_ _27073_/Q _27105_/Q _23845_/S vssd1 vssd1 vccd1 vccd1 _23830_/X sky130_fd_sc_hd__mux2_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater342 _27756_/CLK vssd1 vssd1 vccd1 vccd1 _27758_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater353 _27577_/CLK vssd1 vssd1 vccd1 vccd1 _27584_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater364 _27377_/CLK vssd1 vssd1 vccd1 vccd1 _27681_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater375 _27454_/CLK vssd1 vssd1 vccd1 vccd1 _27458_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater386 _27353_/CLK vssd1 vssd1 vccd1 vccd1 _27105_/CLK sky130_fd_sc_hd__clkbuf_1
X_23761_ _23860_/A vssd1 vssd1 vccd1 vccd1 _23761_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater397 _27443_/CLK vssd1 vssd1 vccd1 vccd1 _27473_/CLK sky130_fd_sc_hd__clkbuf_1
X_20973_ _21145_/A vssd1 vssd1 vccd1 vccd1 _21040_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25500_ _25560_/A vssd1 vssd1 vccd1 vccd1 _25500_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22712_ _22712_/A vssd1 vssd1 vccd1 vccd1 _22712_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26480_ _20998_/X _26480_/D vssd1 vssd1 vccd1 vccd1 _26480_/Q sky130_fd_sc_hd__dfxtp_1
X_23692_ _24906_/A _27251_/Q _23694_/S vssd1 vssd1 vccd1 vccd1 _23693_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25431_ _25474_/A vssd1 vssd1 vccd1 vccd1 _25431_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22643_ _22630_/X _22632_/X _22634_/X _22636_/X _22637_/X _22638_/X vssd1 vssd1 vccd1
+ vccd1 _22644_/A sky130_fd_sc_hd__mux4_1
XFILLER_90_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25362_ _25362_/A vssd1 vssd1 vccd1 vccd1 _27721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22574_ _22574_/A vssd1 vssd1 vccd1 vccd1 _22574_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24313_ _27541_/Q _24317_/B vssd1 vssd1 vccd1 vccd1 _24314_/A sky130_fd_sc_hd__and2_1
X_27101_ _27415_/CLK _27101_/D vssd1 vssd1 vccd1 vccd1 _27101_/Q sky130_fd_sc_hd__dfxtp_1
X_21525_ _21513_/X _21514_/X _21515_/X _21516_/X _21517_/X _21518_/X vssd1 vssd1 vccd1
+ vccd1 _21526_/A sky130_fd_sc_hd__mux4_1
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25293_ _25323_/A _27510_/Q vssd1 vssd1 vccd1 vccd1 _25295_/A sky130_fd_sc_hd__xor2_2
XFILLER_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27032_ _22918_/X _27032_/D vssd1 vssd1 vccd1 vccd1 _27032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24244_ _24244_/A vssd1 vssd1 vccd1 vccd1 _27393_/D sky130_fd_sc_hd__clkbuf_1
X_21456_ _21456_/A vssd1 vssd1 vccd1 vccd1 _21456_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20407_ _20407_/A vssd1 vssd1 vccd1 vccd1 _20407_/X sky130_fd_sc_hd__clkbuf_1
X_24175_ _24175_/A vssd1 vssd1 vccd1 vccd1 _24184_/B sky130_fd_sc_hd__clkbuf_1
X_21387_ _21373_/X _21374_/X _21375_/X _21376_/X _21377_/X _21378_/X vssd1 vssd1 vccd1
+ vccd1 _21388_/A sky130_fd_sc_hd__mux4_1
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23126_ _27104_/Q _17696_/X _23132_/S vssd1 vssd1 vccd1 vccd1 _23127_/A sky130_fd_sc_hd__mux2_1
X_20338_ _20338_/A vssd1 vssd1 vccd1 vccd1 _20412_/A sky130_fd_sc_hd__buf_2
X_27934_ _27934_/A _15949_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_23057_ _27074_/Q _17702_/X _23059_/S vssd1 vssd1 vccd1 vccd1 _23058_/A sky130_fd_sc_hd__mux2_1
X_20269_ _20335_/A vssd1 vssd1 vccd1 vccd1 _20269_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22008_ _22008_/A vssd1 vssd1 vccd1 vccd1 _22008_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26816_ _22166_/X _26816_/D vssd1 vssd1 vccd1 vccd1 _26816_/Q sky130_fd_sc_hd__dfxtp_1
X_14830_ _14830_/A vssd1 vssd1 vccd1 vccd1 _26515_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27796_ _25634_/X _27796_/D vssd1 vssd1 vccd1 vccd1 _27796_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26747_ _21924_/X _26747_/D vssd1 vssd1 vccd1 vccd1 _26747_/Q sky130_fd_sc_hd__dfxtp_1
X_14761_ _14759_/X _26538_/Q _14773_/S vssd1 vssd1 vccd1 vccd1 _14762_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23959_ _23943_/X _23953_/X _23957_/X _23958_/X vssd1 vssd1 vccd1 vccd1 _27291_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16500_ _16500_/A _16500_/B vssd1 vssd1 vccd1 vccd1 _16700_/B sky130_fd_sc_hd__nor2_1
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _26893_/Q _13710_/X _13705_/X _13711_/Y vssd1 vssd1 vccd1 vccd1 _26893_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ _17479_/X _25828_/Q _17486_/S vssd1 vssd1 vccd1 vccd1 _17481_/A sky130_fd_sc_hd__mux2_1
X_14692_ _26561_/Q _14685_/X _14679_/X _14691_/Y vssd1 vssd1 vccd1 vccd1 _26561_/D
+ sky130_fd_sc_hd__a31o_1
X_26678_ _21686_/X _26678_/D vssd1 vssd1 vccd1 vccd1 _26678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16431_ _16786_/B _16476_/B vssd1 vssd1 vccd1 vccd1 _16719_/C sky130_fd_sc_hd__xnor2_1
XFILLER_108_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13643_ _13913_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13643_/Y sky130_fd_sc_hd__nor2_1
X_25629_ _23025_/X _23026_/X _23027_/X _23028_/X _23029_/X _23030_/X vssd1 vssd1 vccd1
+ vccd1 _25630_/A sky130_fd_sc_hd__mux4_1
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19150_ _19147_/X _19149_/X _19173_/S vssd1 vssd1 vccd1 vccd1 _19150_/X sky130_fd_sc_hd__mux2_1
X_13574_ _26940_/Q _13558_/X _13553_/X _13573_/Y vssd1 vssd1 vccd1 vccd1 _26940_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _16395_/A _16395_/B vssd1 vssd1 vccd1 vccd1 _16851_/A sky130_fd_sc_hd__and2_1
XFILLER_158_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18101_ _18403_/A vssd1 vssd1 vccd1 vccd1 _18101_/X sky130_fd_sc_hd__buf_2
XFILLER_40_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _26307_/Q _13392_/X _15317_/S vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__mux2_1
X_16293_ _27402_/Q _16144_/B _16138_/Y _13085_/A vssd1 vssd1 vccd1 vccd1 _16293_/X
+ sky130_fd_sc_hd__a22o_1
X_19081_ _19078_/X _19079_/X _19173_/S vssd1 vssd1 vccd1 vccd1 _19081_/X sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18032_ _26945_/Q _26913_/Q _26881_/Q _26849_/Q _17922_/X _17951_/X vssd1 vssd1 vccd1
+ vccd1 _18032_/X sky130_fd_sc_hd__mux4_2
XFILLER_200_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15244_ _15244_/A vssd1 vssd1 vccd1 vccd1 _26338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15175_ _15175_/A vssd1 vssd1 vccd1 vccd1 _15184_/S sky130_fd_sc_hd__clkbuf_2
X_14126_ _26755_/Q _14117_/X _14120_/X _14125_/Y vssd1 vssd1 vccd1 vccd1 _26755_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19983_ _19983_/A vssd1 vssd1 vccd1 vccd1 _19983_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14057_ _26779_/Q _14042_/X _13954_/B _14056_/Y vssd1 vssd1 vccd1 vccd1 _26779_/D
+ sky130_fd_sc_hd__a31o_1
X_18934_ _18801_/X _18925_/X _18928_/X _18933_/X _18840_/X vssd1 vssd1 vccd1 vccd1
+ _18935_/C sky130_fd_sc_hd__a221o_1
XFILLER_140_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13008_ _13008_/A vssd1 vssd1 vccd1 vccd1 _27795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18865_ _18862_/X _18864_/X _19539_/S vssd1 vssd1 vccd1 vccd1 _18865_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17816_ _18384_/A vssd1 vssd1 vccd1 vccd1 _24394_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_11_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18796_ _27793_/Q _26554_/Q _26426_/Q _26106_/Q _18793_/X _18795_/X vssd1 vssd1 vccd1
+ vccd1 _18796_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17747_ _27430_/Q vssd1 vssd1 vccd1 vccd1 _17747_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14959_ _14975_/A vssd1 vssd1 vccd1 vccd1 _15043_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17678_ _25912_/Q _17673_/X _17690_/S vssd1 vssd1 vccd1 vccd1 _17679_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19417_ _19409_/X _19411_/X _19416_/X _19324_/X _19393_/X vssd1 vssd1 vccd1 vccd1
+ _19426_/B sky130_fd_sc_hd__a221o_1
X_16629_ _16666_/B _16629_/B vssd1 vssd1 vccd1 vccd1 _16629_/X sky130_fd_sc_hd__and2_1
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19348_ _19482_/A vssd1 vssd1 vccd1 vccd1 _19348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19279_ _19272_/X _19275_/X _19278_/X _19186_/X _19258_/X vssd1 vssd1 vccd1 vccd1
+ _19292_/B sky130_fd_sc_hd__a221o_1
XFILLER_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21310_ _21378_/A vssd1 vssd1 vccd1 vccd1 _21310_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22290_ _22290_/A vssd1 vssd1 vccd1 vccd1 _22290_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21241_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21241_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21172_ _21172_/A vssd1 vssd1 vccd1 vccd1 _21172_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20123_ _20123_/A vssd1 vssd1 vccd1 vccd1 _20123_/X sky130_fd_sc_hd__clkbuf_1
X_25980_ _25980_/CLK _25980_/D vssd1 vssd1 vccd1 vccd1 _25980_/Q sky130_fd_sc_hd__dfxtp_1
X_20054_ _20044_/X _20045_/X _20046_/X _20047_/X _20048_/X _20049_/X vssd1 vssd1 vccd1
+ vccd1 _20055_/A sky130_fd_sc_hd__mux4_1
X_24931_ _27776_/Q _24931_/B vssd1 vssd1 vccd1 vccd1 _24932_/B sky130_fd_sc_hd__nor2_1
XFILLER_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27650_ _27659_/CLK _27650_/D vssd1 vssd1 vccd1 vccd1 _27650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24862_ _24862_/A _24867_/C vssd1 vssd1 vccd1 vccd1 _24863_/B sky130_fd_sc_hd__xnor2_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater150 _27791_/CLK vssd1 vssd1 vccd1 vccd1 _27420_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26601_ _21420_/X _26601_/D vssd1 vssd1 vccd1 vccd1 _26601_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater161 _27133_/CLK vssd1 vssd1 vccd1 vccd1 _27407_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater172 _27142_/CLK vssd1 vssd1 vccd1 vccd1 _27840_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23813_ _23861_/A vssd1 vssd1 vccd1 vccd1 _23813_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24793_ _27630_/Q _24785_/X _24792_/Y _24787_/X vssd1 vssd1 vccd1 vccd1 _27630_/D
+ sky130_fd_sc_hd__o211a_1
X_27581_ _27642_/CLK _27581_/D vssd1 vssd1 vccd1 vccd1 _27581_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater183 _27832_/CLK vssd1 vssd1 vccd1 vccd1 _27135_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater194 _26017_/CLK vssd1 vssd1 vccd1 vccd1 _25985_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_206 _14503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _14524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23744_ _23744_/A vssd1 vssd1 vccd1 vccd1 _23744_/X sky130_fd_sc_hd__clkbuf_2
X_26532_ _21174_/X _26532_/D vssd1 vssd1 vccd1 vccd1 _26532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _24511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20956_ _20956_/A vssd1 vssd1 vccd1 vccd1 _20956_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_239 _17376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23675_ _27763_/Q _27243_/Q _23683_/S vssd1 vssd1 vccd1 vccd1 _23676_/A sky130_fd_sc_hd__mux2_1
X_26463_ _20934_/X _26463_/D vssd1 vssd1 vccd1 vccd1 _26463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _21145_/A vssd1 vssd1 vccd1 vccd1 _20954_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22626_ _22626_/A vssd1 vssd1 vccd1 vccd1 _22626_/X sky130_fd_sc_hd__clkbuf_1
X_25414_ _25414_/A vssd1 vssd1 vccd1 vccd1 _27745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26394_ _20683_/X _26394_/D vssd1 vssd1 vccd1 vccd1 _26394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25345_ _27718_/Q _25308_/X _25344_/Y _13423_/X vssd1 vssd1 vccd1 vccd1 _27718_/D
+ sky130_fd_sc_hd__o211a_1
X_22557_ _22539_/X _22542_/X _22545_/X _22548_/X _22549_/X _22550_/X vssd1 vssd1 vccd1
+ vccd1 _22558_/A sky130_fd_sc_hd__mux4_1
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21508_ _21508_/A vssd1 vssd1 vccd1 vccd1 _21508_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25276_ _25323_/A _27508_/Q vssd1 vssd1 vccd1 vccd1 _25282_/A sky130_fd_sc_hd__xor2_2
X_13290_ _13290_/A vssd1 vssd1 vccd1 vccd1 _27015_/D sky130_fd_sc_hd__clkbuf_1
X_22488_ _22520_/A vssd1 vssd1 vccd1 vccd1 _22488_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27015_ _22860_/X _27015_/D vssd1 vssd1 vccd1 vccd1 _27015_/Q sky130_fd_sc_hd__dfxtp_1
X_24227_ _24227_/A vssd1 vssd1 vccd1 vccd1 _27383_/D sky130_fd_sc_hd__clkbuf_1
X_21439_ _21427_/X _21428_/X _21429_/X _21430_/X _21431_/X _21432_/X vssd1 vssd1 vccd1
+ vccd1 _21440_/A sky130_fd_sc_hd__mux4_1
XFILLER_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24158_ _27456_/Q _24162_/B vssd1 vssd1 vccd1 vccd1 _24159_/A sky130_fd_sc_hd__and2_1
XFILLER_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23109_ _23109_/A _25735_/B _23109_/C vssd1 vssd1 vccd1 vccd1 _24002_/A sky130_fd_sc_hd__and3_2
X_24089_ _27393_/Q _24095_/B vssd1 vssd1 vccd1 vccd1 _24090_/A sky130_fd_sc_hd__and2_1
XFILLER_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16980_ _24624_/B _16982_/C _16980_/C vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__and3_1
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ input1/X vssd1 vssd1 vccd1 vccd1 _15956_/A sky130_fd_sc_hd__clkbuf_4
X_27917_ _27917_/A _15973_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18650_ _25991_/Q _17718_/X _18652_/S vssd1 vssd1 vccd1 vccd1 _18651_/A sky130_fd_sc_hd__mux2_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27848_ _27849_/CLK _27848_/D vssd1 vssd1 vccd1 vccd1 _27848_/Q sky130_fd_sc_hd__dfxtp_1
X_15862_ _15862_/A vssd1 vssd1 vccd1 vccd1 _15862_/Y sky130_fd_sc_hd__inv_2
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ _24061_/A _27380_/Q _17601_/C vssd1 vssd1 vccd1 vccd1 _17658_/A sky130_fd_sc_hd__or3_4
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14813_ _14885_/A _14813_/B vssd1 vssd1 vccd1 vccd1 _14870_/A sky130_fd_sc_hd__nor2_2
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18581_ _18575_/X _18577_/X _18580_/X _18150_/A _18238_/A vssd1 vssd1 vccd1 vccd1
+ _18582_/C sky130_fd_sc_hd__a221o_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27779_ _27781_/CLK _27779_/D vssd1 vssd1 vccd1 vccd1 _27779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15793_ _15793_/A vssd1 vssd1 vccd1 vccd1 _26102_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17532_ _17408_/X _25843_/Q _17540_/S vssd1 vssd1 vccd1 vccd1 _17533_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _14811_/S vssd1 vssd1 vccd1 vccd1 _14757_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17463_ _27420_/Q vssd1 vssd1 vccd1 vccd1 _17463_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14675_ _15749_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14675_/Y sky130_fd_sc_hd__nor2_1
X_19202_ _19202_/A vssd1 vssd1 vccd1 vccd1 _26056_/D sky130_fd_sc_hd__clkbuf_1
X_16414_ _25952_/Q _16412_/X _16413_/X vssd1 vssd1 vccd1 vccd1 _16734_/B sky130_fd_sc_hd__a21oi_1
X_13626_ _13639_/A vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17394_ _25655_/A vssd1 vssd1 vccd1 vccd1 _19832_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19133_ _27805_/Q _26566_/Q _26438_/Q _26118_/Q _18922_/X _18901_/X vssd1 vssd1 vccd1
+ vccd1 _19133_/X sky130_fd_sc_hd__mux4_2
Xrepeater75 _27435_/CLK vssd1 vssd1 vccd1 vccd1 _25897_/CLK sky130_fd_sc_hd__clkbuf_1
X_16345_ _16345_/A _16345_/B vssd1 vssd1 vccd1 vccd1 _16347_/B sky130_fd_sc_hd__xnor2_1
XFILLER_157_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater86 _27293_/CLK vssd1 vssd1 vccd1 vccd1 _27296_/CLK sky130_fd_sc_hd__clkbuf_1
X_13557_ _26944_/Q _13535_/X _13553_/X _13556_/Y vssd1 vssd1 vccd1 vccd1 _26944_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_201_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater97 _27121_/CLK vssd1 vssd1 vccd1 vccd1 _26030_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19064_ _19062_/X _19063_/X _19499_/S vssd1 vssd1 vccd1 vccd1 _19064_/X sky130_fd_sc_hd__mux2_1
X_16276_ _16508_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16276_/Y sky130_fd_sc_hd__nor2_1
X_13488_ _27355_/Q _13108_/A _13102_/A _27323_/Q _13120_/X vssd1 vssd1 vccd1 vccd1
+ _16536_/A sky130_fd_sc_hd__a221oi_4
XFILLER_173_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18015_ _18009_/X _18013_/X _18014_/X vssd1 vssd1 vccd1 vccd1 _18015_/X sky130_fd_sc_hd__o21a_1
X_15227_ _15227_/A vssd1 vssd1 vccd1 vccd1 _26346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ _26376_/Q _13376_/X _15162_/S vssd1 vssd1 vccd1 vccd1 _15159_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _26762_/Q _14104_/X _14107_/X _14108_/Y vssd1 vssd1 vccd1 vccd1 _26762_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15089_ _15089_/A vssd1 vssd1 vccd1 vccd1 _26407_/D sky130_fd_sc_hd__clkbuf_1
X_19966_ _19956_/X _19957_/X _19958_/X _19959_/X _19960_/X _19961_/X vssd1 vssd1 vccd1
+ vccd1 _19967_/A sky130_fd_sc_hd__mux4_1
XFILLER_141_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18917_ _18932_/A vssd1 vssd1 vccd1 vccd1 _24405_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_122_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19897_ _19897_/A vssd1 vssd1 vccd1 vccd1 _19897_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18848_ _26683_/Q _26651_/Q _26619_/Q _26587_/Q _18847_/X _18782_/X vssd1 vssd1 vccd1
+ vccd1 _18848_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18779_ _27599_/Q vssd1 vssd1 vccd1 vccd1 _18897_/A sky130_fd_sc_hd__buf_2
XFILLER_36_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20810_ _20791_/X _20795_/X _20799_/X _20803_/X _20804_/X _20805_/X vssd1 vssd1 vccd1
+ vccd1 _20811_/A sky130_fd_sc_hd__mux4_1
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21790_ _21790_/A vssd1 vssd1 vccd1 vccd1 _21790_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20741_ _20773_/A vssd1 vssd1 vccd1 vccd1 _20741_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23460_ _23598_/A vssd1 vssd1 vccd1 vccd1 _25132_/A sky130_fd_sc_hd__clkbuf_2
X_20672_ _20672_/A vssd1 vssd1 vccd1 vccd1 _20672_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22411_ _22401_/X _22402_/X _22403_/X _22404_/X _22405_/X _22406_/X vssd1 vssd1 vccd1
+ vccd1 _22412_/A sky130_fd_sc_hd__mux4_1
XFILLER_32_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23391_ _24790_/A _27254_/Q _27250_/Q _24778_/A vssd1 vssd1 vccd1 vccd1 _23391_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25130_ _25130_/A _25130_/B vssd1 vssd1 vccd1 vccd1 _25131_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22342_ _22342_/A vssd1 vssd1 vccd1 vccd1 _22342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25061_ _27229_/Q vssd1 vssd1 vccd1 vccd1 _25061_/X sky130_fd_sc_hd__buf_2
X_22273_ _22261_/X _22262_/X _22263_/X _22264_/X _22266_/X _22268_/X vssd1 vssd1 vccd1
+ vccd1 _22274_/A sky130_fd_sc_hd__mux4_1
XFILLER_191_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_818 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24012_ _27092_/Q _24001_/X _24002_/X _27124_/Q _24003_/X vssd1 vssd1 vccd1 vccd1
+ _24012_/X sky130_fd_sc_hd__a221o_1
XFILLER_89_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21224_ _21224_/A vssd1 vssd1 vccd1 vccd1 _21224_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21155_ _21144_/X _21146_/X _21148_/X _21150_/X _21151_/X _21152_/X vssd1 vssd1 vccd1
+ vccd1 _21156_/A sky130_fd_sc_hd__mux4_1
XFILLER_144_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20106_ _20095_/X _20097_/X _20099_/X _20101_/X _20102_/X _20103_/X vssd1 vssd1 vccd1
+ vccd1 _20107_/A sky130_fd_sc_hd__mux4_1
X_25963_ _25963_/CLK _25963_/D vssd1 vssd1 vccd1 vccd1 _25963_/Q sky130_fd_sc_hd__dfxtp_1
X_21086_ _21086_/A vssd1 vssd1 vccd1 vccd1 _21086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27702_ _27703_/CLK _27702_/D vssd1 vssd1 vccd1 vccd1 _27702_/Q sky130_fd_sc_hd__dfxtp_1
X_24914_ _24914_/A vssd1 vssd1 vccd1 vccd1 _24914_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20037_ _20037_/A vssd1 vssd1 vccd1 vccd1 _20037_/X sky130_fd_sc_hd__clkbuf_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25894_ _26007_/CLK _25894_/D vssd1 vssd1 vccd1 vccd1 _25894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27633_ _27633_/CLK _27633_/D vssd1 vssd1 vccd1 vccd1 _27633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24845_ _24851_/C _24845_/B vssd1 vssd1 vccd1 vccd1 _24846_/B sky130_fd_sc_hd__or2_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27564_ _27564_/CLK _27564_/D vssd1 vssd1 vccd1 vccd1 _27564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _21988_/A vssd1 vssd1 vccd1 vccd1 _21988_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24776_ _24776_/A _24786_/B vssd1 vssd1 vccd1 vccd1 _24776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26515_ _21116_/X _26515_/D vssd1 vssd1 vccd1 vccd1 _26515_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20939_ _20955_/A vssd1 vssd1 vccd1 vccd1 _20939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23727_ _27370_/Q _24005_/A vssd1 vssd1 vccd1 vccd1 _23728_/A sky130_fd_sc_hd__and2_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27495_ _27495_/CLK _27495_/D vssd1 vssd1 vccd1 vccd1 _27495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14460_ _14530_/A vssd1 vssd1 vccd1 vccd1 _14460_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26446_ _20878_/X _26446_/D vssd1 vssd1 vccd1 vccd1 _26446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23658_ _23658_/A vssd1 vssd1 vccd1 vccd1 _27235_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ _14801_/A vssd1 vssd1 vccd1 vccd1 _13411_/X sky130_fd_sc_hd__buf_4
X_14391_ _26659_/Q _14379_/X _14385_/X _14390_/Y vssd1 vssd1 vccd1 vccd1 _26659_/D
+ sky130_fd_sc_hd__a31o_1
X_22609_ _22609_/A vssd1 vssd1 vccd1 vccd1 _22609_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23589_ _23596_/A _23589_/B vssd1 vssd1 vccd1 vccd1 _23590_/A sky130_fd_sc_hd__and2_1
X_26377_ _20631_/X _26377_/D vssd1 vssd1 vccd1 vccd1 _26377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16130_ _16792_/A vssd1 vssd1 vccd1 vccd1 _16836_/A sky130_fd_sc_hd__clkbuf_2
X_13342_ _26995_/Q _13341_/X _13351_/S vssd1 vssd1 vccd1 vccd1 _13343_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25328_ _25328_/A _25325_/A vssd1 vssd1 vccd1 vccd1 _25329_/D sky130_fd_sc_hd__or2b_1
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_623 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13273_ _13273_/A vssd1 vssd1 vccd1 vccd1 _27023_/D sky130_fd_sc_hd__clkbuf_1
X_16061_ _16056_/Y _27267_/Q _16059_/X _16060_/Y _27265_/Q vssd1 vssd1 vccd1 vccd1
+ _16063_/C sky130_fd_sc_hd__o221a_1
X_25259_ _25249_/A _25252_/B _25267_/A vssd1 vssd1 vccd1 vccd1 _25260_/B sky130_fd_sc_hd__a21bo_1
XFILLER_183_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ _26439_/Q _15002_/X _15003_/X _15011_/Y vssd1 vssd1 vccd1 vccd1 _26439_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_521 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ _19812_/X _19813_/X _19814_/X _19815_/X _19817_/X _19819_/X vssd1 vssd1 vccd1
+ vccd1 _19821_/A sky130_fd_sc_hd__mux4_1
XFILLER_190_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19751_ _19815_/A vssd1 vssd1 vccd1 vccd1 _19751_/X sky130_fd_sc_hd__clkbuf_1
X_16963_ _16971_/B _16979_/B _27592_/Q vssd1 vssd1 vccd1 vccd1 _16963_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18702_ _26014_/Q _17689_/X _18702_/S vssd1 vssd1 vccd1 vccd1 _18703_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15914_ _15918_/A vssd1 vssd1 vccd1 vccd1 _15914_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_652 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19682_ _19714_/A vssd1 vssd1 vccd1 vccd1 _19682_/X sky130_fd_sc_hd__clkbuf_2
X_16894_ _16877_/A _16890_/X _16891_/Y _16893_/Y vssd1 vssd1 vccd1 vccd1 _24232_/A
+ sky130_fd_sc_hd__o31a_1
X_18633_ _25983_/Q _17692_/X _18641_/S vssd1 vssd1 vccd1 vccd1 _18634_/A sky130_fd_sc_hd__mux2_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15845_ _13216_/X _26078_/Q _15849_/S vssd1 vssd1 vccd1 vccd1 _15846_/A sky130_fd_sc_hd__mux2_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ _18842_/A _18564_/B _18564_/C vssd1 vssd1 vccd1 vccd1 _18565_/A sky130_fd_sc_hd__and3_1
XFILLER_80_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _26109_/Q _15774_/X _15766_/X _15775_/Y vssd1 vssd1 vccd1 vccd1 _26109_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12988_/A vssd1 vssd1 vccd1 vccd1 _27804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17515_ _17514_/X _25839_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17516_/A sky130_fd_sc_hd__mux2_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ _14727_/A vssd1 vssd1 vccd1 vccd1 _14727_/X sky130_fd_sc_hd__clkbuf_4
X_18495_ _18493_/X _18494_/X _18532_/S vssd1 vssd1 vccd1 vccd1 _18495_/X sky130_fd_sc_hd__mux2_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17446_ _17446_/A vssd1 vssd1 vccd1 vccd1 _25817_/D sky130_fd_sc_hd__clkbuf_1
X_14658_ _14671_/A vssd1 vssd1 vccd1 vccd1 _14658_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ _26930_/Q _13599_/X _13603_/X _13608_/Y vssd1 vssd1 vccd1 vccd1 _26930_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17377_ _27225_/Q _17376_/X _17387_/S vssd1 vssd1 vccd1 vccd1 _17378_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14589_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14589_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19116_ _19412_/A vssd1 vssd1 vccd1 vccd1 _19116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16328_ _16345_/A vssd1 vssd1 vccd1 vccd1 _16862_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19047_ _19045_/X _19046_/X _19047_/S vssd1 vssd1 vccd1 vccd1 _19047_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16259_ _16502_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19949_ _19949_/A vssd1 vssd1 vccd1 vccd1 _19949_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22960_ _23029_/A vssd1 vssd1 vccd1 vccd1 _22960_/X sky130_fd_sc_hd__clkbuf_2
X_21911_ _21911_/A vssd1 vssd1 vccd1 vccd1 _21911_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22891_ _22891_/A vssd1 vssd1 vccd1 vccd1 _22957_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21842_ _21842_/A vssd1 vssd1 vccd1 vccd1 _21842_/X sky130_fd_sc_hd__clkbuf_1
X_24630_ _24630_/A vssd1 vssd1 vccd1 vccd1 _27573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24561_ _27642_/Q _24565_/B vssd1 vssd1 vccd1 vccd1 _24562_/A sky130_fd_sc_hd__and2_1
X_21773_ _21758_/X _21760_/X _21762_/X _21764_/X _21765_/X _21766_/X vssd1 vssd1 vccd1
+ vccd1 _21774_/A sky130_fd_sc_hd__mux4_1
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26300_ _20367_/X _26300_/D vssd1 vssd1 vccd1 vccd1 _26300_/Q sky130_fd_sc_hd__dfxtp_1
X_20724_ _20772_/A vssd1 vssd1 vccd1 vccd1 _20724_/X sky130_fd_sc_hd__clkbuf_1
X_23512_ _23512_/A vssd1 vssd1 vccd1 vccd1 _27195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24492_ _24551_/S vssd1 vssd1 vccd1 vccd1 _24492_/Y sky130_fd_sc_hd__inv_2
X_27280_ _27379_/CLK _27280_/D vssd1 vssd1 vccd1 vccd1 _27280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23443_ _27171_/Q _23443_/B vssd1 vssd1 vccd1 vccd1 _23443_/X sky130_fd_sc_hd__or2_1
X_26231_ _20123_/X _26231_/D vssd1 vssd1 vccd1 vccd1 _26231_/Q sky130_fd_sc_hd__dfxtp_1
X_20655_ _20687_/A vssd1 vssd1 vccd1 vccd1 _20655_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23374_ _24947_/A _23363_/Y _23368_/X _23373_/X vssd1 vssd1 vccd1 vccd1 _23374_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_20_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26162_ _19877_/X _26162_/D vssd1 vssd1 vccd1 vccd1 _26162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20586_ _20586_/A vssd1 vssd1 vccd1 vccd1 _20586_/X sky130_fd_sc_hd__buf_2
XFILLER_99_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22325_ _22315_/X _22316_/X _22317_/X _22318_/X _22319_/X _22320_/X vssd1 vssd1 vccd1
+ vccd1 _22326_/A sky130_fd_sc_hd__mux4_1
XFILLER_125_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25113_ _25113_/A _25356_/A vssd1 vssd1 vccd1 vccd1 _25113_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26093_ _19634_/X _26093_/D vssd1 vssd1 vccd1 vccd1 _26093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25044_ _27834_/Q _27138_/Q _25883_/Q _25851_/Q _25018_/X _25035_/X vssd1 vssd1 vccd1
+ vccd1 _25044_/X sky130_fd_sc_hd__mux4_1
X_22256_ _22256_/A vssd1 vssd1 vccd1 vccd1 _22256_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21207_ _21195_/X _21196_/X _21197_/X _21198_/X _21199_/X _21200_/X vssd1 vssd1 vccd1
+ vccd1 _21208_/A sky130_fd_sc_hd__mux4_1
XFILLER_151_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22187_ _22173_/X _22174_/X _22175_/X _22176_/X _22179_/X _22182_/X vssd1 vssd1 vccd1
+ vccd1 _22188_/A sky130_fd_sc_hd__mux4_1
XFILLER_160_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21138_ _21138_/A vssd1 vssd1 vccd1 vccd1 _21138_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26995_ _22792_/X _26995_/D vssd1 vssd1 vccd1 vccd1 _26995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13960_ _26806_/Q _13949_/X _13944_/X _13959_/Y vssd1 vssd1 vccd1 vccd1 _26806_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21069_ _21058_/X _21060_/X _21062_/X _21064_/X _21065_/X _21066_/X vssd1 vssd1 vccd1
+ vccd1 _21070_/A sky130_fd_sc_hd__mux4_1
X_25946_ _27356_/CLK _25946_/D vssd1 vssd1 vccd1 vccd1 _25946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13891_ _13891_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13891_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25877_ _27133_/CLK _25877_/D vssd1 vssd1 vccd1 vccd1 _25877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27616_ _27617_/CLK _27616_/D vssd1 vssd1 vccd1 vccd1 _27616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ _13067_/X _26167_/Q _15634_/S vssd1 vssd1 vccd1 vccd1 _15631_/A sky130_fd_sc_hd__mux2_1
X_24828_ _24828_/A _24828_/B _24828_/C vssd1 vssd1 vccd1 vccd1 _24829_/A sky130_fd_sc_hd__and3_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27547_ _27564_/CLK _27547_/D vssd1 vssd1 vccd1 vccd1 _27547_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15561_/A vssd1 vssd1 vccd1 vccd1 _26198_/D sky130_fd_sc_hd__clkbuf_1
X_24759_ _24759_/A _24759_/B vssd1 vssd1 vccd1 vccd1 _24759_/Y sky130_fd_sc_hd__nand2_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _27850_/Q _27154_/Q _25899_/Q _25867_/Q _17264_/X _17252_/X vssd1 vssd1 vccd1
+ vccd1 _17300_/X sky130_fd_sc_hd__mux4_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _15767_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14512_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18280_ _26283_/Q _26251_/Q _26219_/Q _26187_/Q _18185_/X _18209_/X vssd1 vssd1 vccd1
+ vccd1 _18280_/X sky130_fd_sc_hd__mux4_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_872 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27478_ _27478_/CLK _27478_/D vssd1 vssd1 vccd1 vccd1 _27478_/Q sky130_fd_sc_hd__dfxtp_1
X_15492_ _15549_/S vssd1 vssd1 vccd1 vccd1 _15501_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _25829_/Q _26028_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17231_/X sky130_fd_sc_hd__mux2_1
X_14443_ _15716_/A _14446_/B vssd1 vssd1 vccd1 vccd1 _14443_/Y sky130_fd_sc_hd__nor2_1
X_26429_ _20815_/X _26429_/D vssd1 vssd1 vccd1 vccd1 _26429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17162_ _27078_/Q _27110_/Q _17173_/S vssd1 vssd1 vccd1 vccd1 _17162_/X sky130_fd_sc_hd__mux2_1
X_14374_ _14374_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14374_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ _16201_/A vssd1 vssd1 vccd1 vccd1 _16191_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13325_ _14715_/A vssd1 vssd1 vccd1 vccd1 _13325_/X sky130_fd_sc_hd__buf_2
XFILLER_183_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17093_ _27833_/Q _27137_/Q _25882_/Q _25850_/Q _17081_/X _17069_/X vssd1 vssd1 vccd1
+ vccd1 _17093_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16044_ _27476_/Q _27372_/Q vssd1 vssd1 vccd1 vccd1 _16044_/X sky130_fd_sc_hd__or2_1
X_13256_ _27030_/Q _13072_/X _13258_/S vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13187_ _27279_/Q _13201_/B vssd1 vssd1 vccd1 vccd1 _13187_/X sky130_fd_sc_hd__and2_1
XFILLER_123_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19803_ _19803_/A vssd1 vssd1 vccd1 vccd1 _19803_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17995_ _18468_/A vssd1 vssd1 vccd1 vccd1 _17995_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19734_ _19726_/X _19727_/X _19728_/X _19729_/X _19731_/X _19733_/X vssd1 vssd1 vccd1
+ vccd1 _19735_/A sky130_fd_sc_hd__mux4_1
X_16946_ _16927_/X _16930_/X _16936_/X _16945_/X vssd1 vssd1 vccd1 vccd1 _16947_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_42_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19665_ _19729_/A vssd1 vssd1 vccd1 vccd1 _19665_/X sky130_fd_sc_hd__clkbuf_1
X_16877_ _16877_/A vssd1 vssd1 vccd1 vccd1 _16877_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18616_ _25977_/Q vssd1 vssd1 vccd1 vccd1 _24825_/A sky130_fd_sc_hd__inv_2
X_27986__452 vssd1 vssd1 vccd1 vccd1 _27986__452/HI _27986_/A sky130_fd_sc_hd__conb_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _15828_/A vssd1 vssd1 vccd1 vccd1 _26086_/D sky130_fd_sc_hd__clkbuf_1
X_19596_ _19596_/A vssd1 vssd1 vccd1 vccd1 _19596_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18547_ _18547_/A vssd1 vssd1 vccd1 vccd1 _25973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15759_ _26115_/Q _15747_/X _15753_/X _15758_/Y vssd1 vssd1 vccd1 vccd1 _26115_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18478_ _26164_/Q _26100_/Q _27028_/Q _26996_/Q _18455_/X _18387_/X vssd1 vssd1 vccd1
+ vccd1 _18480_/A sky130_fd_sc_hd__mux4_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17429_ _17428_/X _25812_/Q _17438_/S vssd1 vssd1 vccd1 vccd1 _17430_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20440_ _20424_/X _20425_/X _20426_/X _20427_/X _20430_/X _20433_/X vssd1 vssd1 vccd1
+ vccd1 _20441_/A sky130_fd_sc_hd__mux4_1
XFILLER_20_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ _20371_/A vssd1 vssd1 vccd1 vccd1 _20371_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22110_ _22546_/A vssd1 vssd1 vccd1 vccd1 _22457_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_23090_ _27089_/Q _17750_/X _23092_/S vssd1 vssd1 vccd1 vccd1 _23091_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22041_ _22035_/X _22036_/X _22037_/X _22038_/X _22039_/X _22040_/X vssd1 vssd1 vccd1
+ vccd1 _22042_/A sky130_fd_sc_hd__mux4_1
XFILLER_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25800_ _25800_/A vssd1 vssd1 vccd1 vccd1 _27854_/D sky130_fd_sc_hd__clkbuf_1
X_26780_ _22042_/X _26780_/D vssd1 vssd1 vccd1 vccd1 _26780_/Q sky130_fd_sc_hd__dfxtp_1
X_23992_ _27851_/Q _27155_/Q _25900_/Q _25868_/Q _23967_/X _23991_/X vssd1 vssd1 vccd1
+ vccd1 _23992_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25731_ _25721_/X _25722_/X _25723_/X _25724_/X _25725_/X _25726_/X vssd1 vssd1 vccd1
+ vccd1 _25732_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22943_ _22943_/A vssd1 vssd1 vccd1 vccd1 _22943_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_997 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25662_ _25710_/A vssd1 vssd1 vccd1 vccd1 _25662_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22874_ _22943_/A vssd1 vssd1 vccd1 vccd1 _22874_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27401_ _27401_/CLK _27401_/D vssd1 vssd1 vccd1 vccd1 _27401_/Q sky130_fd_sc_hd__dfxtp_1
X_24613_ _24613_/A vssd1 vssd1 vccd1 vccd1 _27565_/D sky130_fd_sc_hd__clkbuf_1
X_21825_ _21825_/A vssd1 vssd1 vccd1 vccd1 _21825_/X sky130_fd_sc_hd__clkbuf_1
X_25593_ _24804_/A _25564_/X _25590_/X _25591_/Y _25592_/X vssd1 vssd1 vccd1 vccd1
+ _27779_/D sky130_fd_sc_hd__a221oi_1
XFILLER_197_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27332_ _27332_/CLK _27332_/D vssd1 vssd1 vccd1 vccd1 _27332_/Q sky130_fd_sc_hd__dfxtp_1
X_21756_ _21756_/A vssd1 vssd1 vccd1 vccd1 _21756_/X sky130_fd_sc_hd__clkbuf_1
X_24544_ _24544_/A vssd1 vssd1 vccd1 vccd1 _27535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20707_ _20772_/A vssd1 vssd1 vccd1 vccd1 _20707_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27263_ _27263_/CLK _27263_/D vssd1 vssd1 vccd1 vccd1 _27263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21687_ _21667_/X _21670_/X _21673_/X _21676_/X _21677_/X _21678_/X vssd1 vssd1 vccd1
+ vccd1 _21688_/A sky130_fd_sc_hd__mux4_1
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24475_ _24475_/A vssd1 vssd1 vccd1 vccd1 _27513_/D sky130_fd_sc_hd__clkbuf_1
X_26214_ _20059_/X _26214_/D vssd1 vssd1 vccd1 vccd1 _26214_/Q sky130_fd_sc_hd__dfxtp_1
X_20638_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20638_/X sky130_fd_sc_hd__clkbuf_1
X_23426_ input31/X _23415_/X _23425_/X _23421_/X vssd1 vssd1 vccd1 vccd1 _27164_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27194_ _27578_/CLK _27194_/D vssd1 vssd1 vccd1 vccd1 _27194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23357_ _27780_/Q vssd1 vssd1 vccd1 vccd1 _24806_/A sky130_fd_sc_hd__inv_2
X_26145_ _19821_/X _26145_/D vssd1 vssd1 vccd1 vccd1 _26145_/Q sky130_fd_sc_hd__dfxtp_1
X_20569_ _20601_/A vssd1 vssd1 vccd1 vccd1 _20569_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22308_ _22308_/A vssd1 vssd1 vccd1 vccd1 _22308_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13110_ _27357_/Q _13108_/X _13029_/A _27325_/Q _13109_/X vssd1 vssd1 vccd1 vccd1
+ _14740_/A sky130_fd_sc_hd__a221o_4
XFILLER_192_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14090_ _14090_/A vssd1 vssd1 vccd1 vccd1 _14090_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23288_ input68/X vssd1 vssd1 vccd1 vccd1 _23288_/Y sky130_fd_sc_hd__inv_2
X_26076_ _19582_/X _26076_/D vssd1 vssd1 vccd1 vccd1 _26076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ _27268_/Q vssd1 vssd1 vccd1 vccd1 _16014_/B sky130_fd_sc_hd__clkbuf_4
X_22239_ _22229_/X _22230_/X _22231_/X _22232_/X _22233_/X _22234_/X vssd1 vssd1 vccd1
+ vccd1 _22240_/A sky130_fd_sc_hd__mux4_1
X_25027_ _27230_/Q vssd1 vssd1 vccd1 vccd1 _25027_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16800_ _16800_/A _16800_/B _16800_/C _16800_/D vssd1 vssd1 vccd1 vccd1 _16812_/A
+ sky130_fd_sc_hd__nor4_1
XFILLER_121_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17780_ _27593_/Q vssd1 vssd1 vccd1 vccd1 _18360_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14992_ _15730_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14992_/Y sky130_fd_sc_hd__nor2_1
X_26978_ _22732_/X _26978_/D vssd1 vssd1 vccd1 vccd1 _26978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16731_ _16731_/A _16731_/B vssd1 vssd1 vccd1 vccd1 _16732_/A sky130_fd_sc_hd__nand2_1
X_25929_ _25995_/CLK _25929_/D vssd1 vssd1 vccd1 vccd1 _25929_/Q sky130_fd_sc_hd__dfxtp_1
X_13943_ _13964_/A vssd1 vssd1 vccd1 vccd1 _14060_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19450_ _19471_/A _19450_/B _19450_/C vssd1 vssd1 vccd1 vccd1 _19451_/A sky130_fd_sc_hd__and3_1
XFILLER_189_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16662_ _16662_/A _16662_/B vssd1 vssd1 vccd1 vccd1 _16662_/X sky130_fd_sc_hd__xor2_1
X_13874_ _13874_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13874_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18401_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18401_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15613_ _26174_/Q _14798_/A _15617_/S vssd1 vssd1 vccd1 vccd1 _15614_/A sky130_fd_sc_hd__mux2_1
X_19381_ _19471_/A _19381_/B _19381_/C vssd1 vssd1 vccd1 vccd1 _19382_/A sky130_fd_sc_hd__and3_1
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16593_ _16593_/A _16593_/B vssd1 vssd1 vccd1 vccd1 _16594_/A sky130_fd_sc_hd__and2_1
X_18332_ _18323_/X _18327_/X _18331_/X _18285_/X _18238_/X vssd1 vssd1 vccd1 vccd1
+ _18333_/C sky130_fd_sc_hd__a221o_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _15544_/A vssd1 vssd1 vccd1 vccd1 _26205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18256_/X _18258_/X _18262_/X _18168_/X _18238_/X vssd1 vssd1 vccd1 vccd1
+ _18264_/C sky130_fd_sc_hd__a221o_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15475_ _26235_/Q _13417_/X _15477_/S vssd1 vssd1 vccd1 vccd1 _15476_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17214_ _17214_/A vssd1 vssd1 vccd1 vccd1 _27932_/A sky130_fd_sc_hd__clkbuf_1
X_14426_ _15703_/A _14426_/B vssd1 vssd1 vccd1 vccd1 _14426_/Y sky130_fd_sc_hd__nor2_1
X_18194_ _18194_/A vssd1 vssd1 vccd1 vccd1 _25957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17145_ _25923_/Q _25989_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17146_/B sky130_fd_sc_hd__mux2_1
X_14357_ _26672_/Q _14352_/X _14345_/X _14356_/Y vssd1 vssd1 vccd1 vccd1 _26672_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_498 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13308_ _13308_/A vssd1 vssd1 vccd1 vccd1 _27007_/D sky130_fd_sc_hd__clkbuf_1
X_17076_ _27071_/Q _27103_/Q _17112_/S vssd1 vssd1 vccd1 vccd1 _17076_/X sky130_fd_sc_hd__mux2_1
X_14288_ _26697_/Q _14283_/X _14284_/X _14287_/Y vssd1 vssd1 vccd1 vccd1 _26697_/D
+ sky130_fd_sc_hd__a31o_1
X_16027_ _16264_/B vssd1 vssd1 vccd1 vccd1 _16287_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13239_ _16182_/A vssd1 vssd1 vccd1 vccd1 _14810_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_522 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17978_ _18156_/A vssd1 vssd1 vccd1 vccd1 _17978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19717_ _19717_/A vssd1 vssd1 vccd1 vccd1 _19717_/X sky130_fd_sc_hd__clkbuf_1
X_16929_ _27487_/Q vssd1 vssd1 vccd1 vccd1 _24209_/A sky130_fd_sc_hd__inv_2
XFILLER_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19648_ _19637_/X _19638_/X _19639_/X _19640_/X _19644_/X _19647_/X vssd1 vssd1 vccd1
+ vccd1 _19649_/A sky130_fd_sc_hd__mux4_1
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19579_ _19570_/X _19572_/X _19574_/X _19576_/X _19577_/X _19578_/X vssd1 vssd1 vccd1
+ vccd1 _19580_/A sky130_fd_sc_hd__mux4_1
XFILLER_81_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21610_ _21610_/A vssd1 vssd1 vccd1 vccd1 _21610_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22590_ _22590_/A vssd1 vssd1 vccd1 vccd1 _22590_/X sky130_fd_sc_hd__clkbuf_1
X_21541_ _21529_/X _21530_/X _21531_/X _21532_/X _21533_/X _21534_/X vssd1 vssd1 vccd1
+ vccd1 _21542_/A sky130_fd_sc_hd__mux4_1
XFILLER_166_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24260_ _24260_/A vssd1 vssd1 vccd1 vccd1 _27402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21472_ _21472_/A vssd1 vssd1 vccd1 vccd1 _21472_/X sky130_fd_sc_hd__clkbuf_1
X_23211_ _17463_/X _27142_/Q _23215_/S vssd1 vssd1 vccd1 vccd1 _23212_/A sky130_fd_sc_hd__mux2_1
X_20423_ _20423_/A vssd1 vssd1 vccd1 vccd1 _20423_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24191_ _27471_/Q _24195_/B vssd1 vssd1 vccd1 vccd1 _24192_/A sky130_fd_sc_hd__and2_1
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23142_ _23142_/A vssd1 vssd1 vccd1 vccd1 _27111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20354_ _20424_/A vssd1 vssd1 vccd1 vccd1 _20354_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23073_ _27081_/Q _17724_/X _23081_/S vssd1 vssd1 vccd1 vccd1 _23074_/A sky130_fd_sc_hd__mux2_1
X_27950_ _27950_/A _15926_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
X_20285_ _20285_/A vssd1 vssd1 vccd1 vccd1 _20285_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22024_ _22072_/A vssd1 vssd1 vccd1 vccd1 _22024_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26901_ _22464_/X _26901_/D vssd1 vssd1 vccd1 vccd1 _26901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26832_ _22224_/X _26832_/D vssd1 vssd1 vccd1 vccd1 _26832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26763_ _21978_/X _26763_/D vssd1 vssd1 vccd1 vccd1 _26763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23975_ _27849_/Q _27153_/Q _25898_/Q _25866_/Q _23967_/X _23944_/X vssd1 vssd1 vccd1
+ vccd1 _23975_/X sky130_fd_sc_hd__mux4_1
XFILLER_186_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25714_ _25714_/A vssd1 vssd1 vccd1 vccd1 _25714_/X sky130_fd_sc_hd__clkbuf_1
X_22926_ _22958_/A vssd1 vssd1 vccd1 vccd1 _22926_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26694_ _21736_/X _26694_/D vssd1 vssd1 vccd1 vccd1 _26694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25645_ _25635_/X _25636_/X _25637_/X _25638_/X _25640_/X _25642_/X vssd1 vssd1 vccd1
+ vccd1 _25646_/A sky130_fd_sc_hd__mux4_1
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22857_ _22857_/A vssd1 vssd1 vccd1 vccd1 _22857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21808_ _21808_/A vssd1 vssd1 vccd1 vccd1 _21808_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _26937_/Q _13580_/X _13587_/X _13589_/Y vssd1 vssd1 vccd1 vccd1 _26937_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25576_ _24794_/A _25564_/X _25574_/X _25575_/Y _25557_/X vssd1 vssd1 vccd1 vccd1
+ _27776_/D sky130_fd_sc_hd__a221oi_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22788_ _22857_/A vssd1 vssd1 vccd1 vccd1 _22788_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27315_ _27334_/CLK _27315_/D vssd1 vssd1 vccd1 vccd1 _27315_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24527_ _24554_/A _27590_/Q _24631_/B vssd1 vssd1 vccd1 vccd1 _24528_/B sky130_fd_sc_hd__mux2_1
X_21739_ _21739_/A vssd1 vssd1 vccd1 vccd1 _21739_/X sky130_fd_sc_hd__clkbuf_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27246_ _27261_/CLK _27246_/D vssd1 vssd1 vccd1 vccd1 _27246_/Q sky130_fd_sc_hd__dfxtp_1
X_15260_ _14810_/X _26330_/Q _15260_/S vssd1 vssd1 vccd1 vccd1 _15261_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24458_ _24480_/A vssd1 vssd1 vccd1 vccd1 _24467_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14211_ _26724_/Q _14199_/X _14207_/X _14210_/Y vssd1 vssd1 vccd1 vccd1 _26724_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23409_ _23409_/A _23409_/B _23409_/C _23408_/X vssd1 vssd1 vccd1 vccd1 _23410_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_177_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27177_ _27180_/CLK _27177_/D vssd1 vssd1 vccd1 vccd1 _27177_/Q sky130_fd_sc_hd__dfxtp_1
X_15191_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15260_/S sky130_fd_sc_hd__buf_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24389_ _24389_/A vssd1 vssd1 vccd1 vccd1 _27475_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 _25854_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ _14157_/A vssd1 vssd1 vccd1 vccd1 _14142_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26128_ _19761_/X _26128_/D vssd1 vssd1 vccd1 vccd1 _26128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14073_ _14127_/A vssd1 vssd1 vccd1 vccd1 _14085_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26059_ _26059_/CLK _26059_/D vssd1 vssd1 vccd1 vccd1 _26059_/Q sky130_fd_sc_hd__dfxtp_1
X_18950_ _19482_/A vssd1 vssd1 vccd1 vccd1 _18950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17901_ _18486_/A vssd1 vssd1 vccd1 vccd1 _17901_/X sky130_fd_sc_hd__buf_4
X_13024_ _13194_/A vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18881_ _18872_/X _18874_/X _18878_/X _18854_/X _18880_/X vssd1 vssd1 vccd1 vccd1
+ _18892_/B sky130_fd_sc_hd__a221o_1
XFILLER_117_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17832_ _18358_/A vssd1 vssd1 vccd1 vccd1 _17832_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17763_ _27435_/Q vssd1 vssd1 vccd1 vccd1 _17763_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14975_ _14975_/A vssd1 vssd1 vccd1 vccd1 _15029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19502_ _26838_/Q _26806_/Q _26774_/Q _26742_/Q _18913_/X _18930_/X vssd1 vssd1 vccd1
+ vccd1 _19502_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16714_ _16641_/A _16710_/X _16713_/Y vssd1 vssd1 vccd1 vccd1 _24230_/A sky130_fd_sc_hd__o21a_1
X_13926_ _13926_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _13926_/Y sky130_fd_sc_hd__nor2_1
X_17694_ _25917_/Q _17692_/X _17706_/S vssd1 vssd1 vccd1 vccd1 _17695_/A sky130_fd_sc_hd__mux2_1
X_19433_ _19431_/X _19432_/X _19387_/X vssd1 vssd1 vccd1 vccd1 _19433_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16645_ _16638_/X _16642_/Y _16644_/Y _16626_/X vssd1 vssd1 vccd1 vccd1 _24259_/A
+ sky130_fd_sc_hd__a22o_1
X_13857_ _13857_/A _13861_/B vssd1 vssd1 vccd1 vccd1 _13857_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19364_ _19473_/A vssd1 vssd1 vccd1 vccd1 _19471_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_62_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16576_ _16576_/A _16576_/B vssd1 vssd1 vccd1 vccd1 _16577_/B sky130_fd_sc_hd__nand2_1
X_13788_ _13882_/A _13799_/B vssd1 vssd1 vccd1 vccd1 _13788_/Y sky130_fd_sc_hd__nor2_1
X_18315_ _26829_/Q _26797_/Q _26765_/Q _26733_/Q _18175_/X _18199_/X vssd1 vssd1 vccd1
+ vccd1 _18315_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15527_ _15527_/A vssd1 vssd1 vccd1 vccd1 _26213_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19295_ _27812_/Q _26573_/Q _26445_/Q _26125_/Q _18913_/A _19445_/A vssd1 vssd1 vccd1
+ vccd1 _19295_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18246_ _18405_/A vssd1 vssd1 vccd1 vccd1 _18378_/S sky130_fd_sc_hd__clkbuf_2
X_15458_ _26243_/Q _13392_/X _15462_/S vssd1 vssd1 vccd1 vccd1 _15459_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14409_ _26652_/Q _14405_/X _14398_/X _14408_/Y vssd1 vssd1 vccd1 vccd1 _26652_/D
+ sky130_fd_sc_hd__a31o_1
X_18177_ _18177_/A vssd1 vssd1 vccd1 vccd1 _18177_/X sky130_fd_sc_hd__buf_2
X_15389_ _15389_/A vssd1 vssd1 vccd1 vccd1 _26274_/D sky130_fd_sc_hd__clkbuf_1
X_17128_ _27204_/Q _17127_/X _17128_/S vssd1 vssd1 vccd1 vccd1 _17129_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17059_ _17057_/X _17058_/X _17033_/X vssd1 vssd1 vccd1 vccd1 _17059_/X sky130_fd_sc_hd__a21bo_1
XFILLER_144_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20070_ _20060_/X _20061_/X _20062_/X _20063_/X _20064_/X _20065_/X vssd1 vssd1 vccd1
+ vccd1 _20071_/A sky130_fd_sc_hd__mux4_1
XFILLER_124_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater310 _27472_/CLK vssd1 vssd1 vccd1 vccd1 _27467_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_135_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater321 _27629_/CLK vssd1 vssd1 vccd1 vccd1 _27511_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater332 _27768_/CLK vssd1 vssd1 vccd1 vccd1 _27774_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater343 _27690_/CLK vssd1 vssd1 vccd1 vccd1 _27756_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater354 _27573_/CLK vssd1 vssd1 vccd1 vccd1 _27577_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater365 _27368_/CLK vssd1 vssd1 vccd1 vccd1 _27377_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater376 _27452_/CLK vssd1 vssd1 vccd1 vccd1 _27454_/CLK sky130_fd_sc_hd__clkbuf_1
X_23760_ _24001_/A vssd1 vssd1 vccd1 vccd1 _23860_/A sky130_fd_sc_hd__buf_2
X_20972_ _21039_/A vssd1 vssd1 vccd1 vccd1 _20972_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater387 _27208_/CLK vssd1 vssd1 vccd1 vccd1 _27353_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater398 _27442_/CLK vssd1 vssd1 vccd1 vccd1 _27443_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22711_ _22697_/X _22698_/X _22699_/X _22700_/X _22702_/X _22704_/X vssd1 vssd1 vccd1
+ vccd1 _22712_/A sky130_fd_sc_hd__mux4_1
XFILLER_198_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23691_ _23691_/A vssd1 vssd1 vccd1 vccd1 _27250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25430_ _25430_/A _25430_/B vssd1 vssd1 vccd1 vccd1 _27754_/D sky130_fd_sc_hd__nor2_1
X_22642_ _22642_/A vssd1 vssd1 vccd1 vccd1 _22642_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22573_ _22561_/X _22562_/X _22563_/X _22564_/X _22565_/X _22566_/X vssd1 vssd1 vccd1
+ vccd1 _22574_/A sky130_fd_sc_hd__mux4_1
X_25361_ _27721_/Q input41/X _25369_/S vssd1 vssd1 vccd1 vccd1 _25362_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27100_ _27677_/CLK _27100_/D vssd1 vssd1 vccd1 vccd1 _27100_/Q sky130_fd_sc_hd__dfxtp_1
X_24312_ _24312_/A vssd1 vssd1 vccd1 vccd1 _27440_/D sky130_fd_sc_hd__clkbuf_1
X_21524_ _21524_/A vssd1 vssd1 vccd1 vccd1 _21524_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25292_ _27711_/Q _25263_/X _25291_/Y _25254_/X vssd1 vssd1 vccd1 vccd1 _27711_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_194_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27031_ _22916_/X _27031_/D vssd1 vssd1 vccd1 vccd1 _27031_/Q sky130_fd_sc_hd__dfxtp_1
X_21455_ _21443_/X _21444_/X _21445_/X _21446_/X _21447_/X _21448_/X vssd1 vssd1 vccd1
+ vccd1 _21456_/A sky130_fd_sc_hd__mux4_1
X_24243_ _24243_/A _24250_/B vssd1 vssd1 vccd1 vccd1 _24244_/A sky130_fd_sc_hd__and2_1
XFILLER_108_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20406_ _20392_/X _20393_/X _20394_/X _20395_/X _20396_/X _20397_/X vssd1 vssd1 vccd1
+ vccd1 _20407_/A sky130_fd_sc_hd__mux4_1
XFILLER_181_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24174_ _24174_/A vssd1 vssd1 vccd1 vccd1 _27358_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_21386_ _21386_/A vssd1 vssd1 vccd1 vccd1 _21386_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20337_ _20337_/A vssd1 vssd1 vccd1 vccd1 _20337_/X sky130_fd_sc_hd__clkbuf_1
X_23125_ _23125_/A vssd1 vssd1 vccd1 vccd1 _27103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27933_ _27933_/A _15952_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
X_23056_ _23056_/A vssd1 vssd1 vccd1 vccd1 _27073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20268_ _20268_/A vssd1 vssd1 vccd1 vccd1 _20335_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22007_ _21997_/X _21998_/X _21999_/X _22000_/X _22002_/X _22004_/X vssd1 vssd1 vccd1
+ vccd1 _22008_/A sky130_fd_sc_hd__mux4_1
XFILLER_62_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20199_ _20199_/A vssd1 vssd1 vccd1 vccd1 _20199_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26815_ _22164_/X _26815_/D vssd1 vssd1 vccd1 vccd1 _26815_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27795_ _25632_/X _27795_/D vssd1 vssd1 vccd1 vccd1 _27795_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26746_ _21922_/X _26746_/D vssd1 vssd1 vccd1 vccd1 _26746_/Q sky130_fd_sc_hd__dfxtp_1
X_14760_ _14792_/A vssd1 vssd1 vccd1 vccd1 _14773_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23958_ _24005_/A vssd1 vssd1 vccd1 vccd1 _23958_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13711_ _13891_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13711_/Y sky130_fd_sc_hd__nor2_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22909_ _22957_/A vssd1 vssd1 vccd1 vccd1 _22909_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26677_ _21684_/X _26677_/D vssd1 vssd1 vccd1 vccd1 _26677_/Q sky130_fd_sc_hd__dfxtp_1
X_14691_ _15764_/A _14699_/B vssd1 vssd1 vccd1 vccd1 _14691_/Y sky130_fd_sc_hd__nor2_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23889_ _27840_/Q _27144_/Q _25889_/Q _25857_/Q _23873_/X _23850_/X vssd1 vssd1 vccd1
+ vccd1 _23889_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16430_ _16722_/A _16430_/B vssd1 vssd1 vccd1 vccd1 _16476_/B sky130_fd_sc_hd__xnor2_1
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13642_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13642_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25628_ _25628_/A vssd1 vssd1 vccd1 vccd1 _25628_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16764_/A _16361_/B vssd1 vssd1 vccd1 vccd1 _16395_/B sky130_fd_sc_hd__xor2_1
XFILLER_188_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13573_ _13936_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13573_/Y sky130_fd_sc_hd__nor2_1
X_25559_ _27710_/Q _25539_/X _25540_/X vssd1 vssd1 vccd1 vccd1 _25559_/Y sky130_fd_sc_hd__a21oi_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18100_ _27803_/Q _26564_/Q _26436_/Q _26116_/Q _18099_/X _17949_/X vssd1 vssd1 vccd1
+ vccd1 _18100_/X sky130_fd_sc_hd__mux4_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15312_/A vssd1 vssd1 vccd1 vccd1 _26308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19080_ _19391_/A vssd1 vssd1 vccd1 vccd1 _19173_/S sky130_fd_sc_hd__clkbuf_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16292_ _16824_/A _16292_/B _16292_/C _16292_/D vssd1 vssd1 vccd1 vccd1 _16301_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _27800_/Q _26561_/Q _26433_/Q _26113_/Q _17920_/X _17949_/X vssd1 vssd1 vccd1
+ vccd1 _18031_/X sky130_fd_sc_hd__mux4_2
X_27229_ _27826_/CLK _27229_/D vssd1 vssd1 vccd1 vccd1 _27229_/Q sky130_fd_sc_hd__dfxtp_1
X_15243_ _14785_/X _26338_/Q _15245_/S vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15174_ _15174_/A vssd1 vssd1 vccd1 vccd1 _26369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _14390_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19982_ _19972_/X _19973_/X _19974_/X _19975_/X _19976_/X _19977_/X vssd1 vssd1 vccd1
+ vccd1 _19983_/A sky130_fd_sc_hd__mux4_1
XFILLER_193_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14056_ _14410_/A _14060_/B vssd1 vssd1 vccd1 vccd1 _14056_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18933_ _18929_/X _18931_/X _18932_/X vssd1 vssd1 vccd1 vccd1 _18933_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _27795_/Q _13009_/B vssd1 vssd1 vccd1 vccd1 _13008_/A sky130_fd_sc_hd__and2_1
X_18864_ _26523_/Q _26491_/Q _26459_/Q _27035_/Q _18829_/X _18863_/X vssd1 vssd1 vccd1
+ vccd1 _18864_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17815_ _27596_/Q vssd1 vssd1 vccd1 vccd1 _18384_/A sky130_fd_sc_hd__buf_2
X_18795_ _19321_/A vssd1 vssd1 vccd1 vccd1 _18795_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28011__477 vssd1 vssd1 vccd1 vccd1 _28011__477/HI _28011_/A sky130_fd_sc_hd__conb_1
X_17746_ _17746_/A vssd1 vssd1 vccd1 vccd1 _25933_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14958_ _15695_/A _15695_/B _15695_/C _15190_/A vssd1 vssd1 vccd1 vccd1 _14975_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13909_ _26823_/Q _13906_/X _13899_/X _13908_/Y vssd1 vssd1 vccd1 vccd1 _26823_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17677_ _17776_/S vssd1 vssd1 vccd1 vccd1 _17690_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14889_ _14889_/A vssd1 vssd1 vccd1 vccd1 _26489_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19416_ _19413_/X _19415_/X _19480_/S vssd1 vssd1 vccd1 vccd1 _19416_/X sky130_fd_sc_hd__mux2_1
X_16628_ _16700_/A _16672_/A _16700_/B _16543_/X vssd1 vssd1 vccd1 vccd1 _16664_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_165_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19347_ _19340_/X _19342_/X _19346_/X _19324_/X _19258_/X vssd1 vssd1 vccd1 vccd1
+ _19362_/B sky130_fd_sc_hd__a221o_1
X_16559_ _16559_/A _16648_/B vssd1 vssd1 vccd1 vccd1 _16561_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19278_ _19276_/X _19277_/X _19346_/S vssd1 vssd1 vccd1 vccd1 _19278_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18229_ _26153_/Q _26089_/Q _27017_/Q _26985_/Q _18182_/X _18228_/X vssd1 vssd1 vccd1
+ vccd1 _18230_/A sky130_fd_sc_hd__mux4_1
XFILLER_191_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21240_ _21304_/A vssd1 vssd1 vccd1 vccd1 _21240_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21171_ _21163_/X _21164_/X _21165_/X _21166_/X _21167_/X _21168_/X vssd1 vssd1 vccd1
+ vccd1 _21172_/A sky130_fd_sc_hd__mux4_1
XFILLER_85_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20122_ _20114_/X _20115_/X _20116_/X _20117_/X _20118_/X _20119_/X vssd1 vssd1 vccd1
+ vccd1 _20123_/A sky130_fd_sc_hd__mux4_1
XFILLER_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20053_ _20053_/A vssd1 vssd1 vccd1 vccd1 _20053_/X sky130_fd_sc_hd__clkbuf_1
X_24930_ _27776_/Q _24931_/B vssd1 vssd1 vccd1 vccd1 _24941_/C sky130_fd_sc_hd__and2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24861_ _24861_/A vssd1 vssd1 vccd1 vccd1 _24861_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater140 _27083_/CLK vssd1 vssd1 vccd1 vccd1 _26026_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26600_ _21418_/X _26600_/D vssd1 vssd1 vccd1 vccd1 _26600_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater151 _27418_/CLK vssd1 vssd1 vccd1 vccd1 _27791_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23812_ _23860_/A vssd1 vssd1 vccd1 vccd1 _23812_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater162 _27132_/CLK vssd1 vssd1 vccd1 vccd1 _27133_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater173 _25925_/CLK vssd1 vssd1 vccd1 vccd1 _27142_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27580_ _27584_/CLK _27580_/D vssd1 vssd1 vccd1 vccd1 _27580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24792_ _24792_/A _24800_/B vssd1 vssd1 vccd1 vccd1 _24792_/Y sky130_fd_sc_hd__nand2_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater184 _25917_/CLK vssd1 vssd1 vccd1 vccd1 _27832_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_207 _14507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater195 _25980_/CLK vssd1 vssd1 vccd1 vccd1 _26017_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_218 _14527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26531_ _21172_/X _26531_/D vssd1 vssd1 vccd1 vccd1 _26531_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23743_ _27786_/Q vssd1 vssd1 vccd1 vccd1 _23744_/A sky130_fd_sc_hd__buf_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _20955_/A vssd1 vssd1 vccd1 vccd1 _20955_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _24511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26462_ _20932_/X _26462_/D vssd1 vssd1 vccd1 vccd1 _26462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23674_ _23720_/S vssd1 vssd1 vccd1 vccd1 _23683_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20886_ _20953_/A vssd1 vssd1 vccd1 vccd1 _20886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25413_ _27745_/Q input57/X _25413_/S vssd1 vssd1 vccd1 vccd1 _25414_/A sky130_fd_sc_hd__mux2_1
X_22625_ _22609_/X _22610_/X _22611_/X _22612_/X _22615_/X _22618_/X vssd1 vssd1 vccd1
+ vccd1 _22626_/A sky130_fd_sc_hd__mux4_1
X_26393_ _20681_/X _26393_/D vssd1 vssd1 vccd1 vccd1 _26393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25344_ _25344_/A _25344_/B vssd1 vssd1 vccd1 vccd1 _25344_/Y sky130_fd_sc_hd__nand2_1
X_22556_ _22556_/A vssd1 vssd1 vccd1 vccd1 _22556_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21507_ _21494_/X _21496_/X _21498_/X _21500_/X _21501_/X _21502_/X vssd1 vssd1 vccd1
+ vccd1 _21508_/A sky130_fd_sc_hd__mux4_1
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25275_ _27709_/Q _25263_/X _25274_/Y _25254_/X vssd1 vssd1 vccd1 vccd1 _27709_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22487_ _22519_/A vssd1 vssd1 vccd1 vccd1 _22487_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27014_ _22852_/X _27014_/D vssd1 vssd1 vccd1 vccd1 _27014_/Q sky130_fd_sc_hd__dfxtp_1
X_24226_ _24226_/A _24233_/B vssd1 vssd1 vccd1 vccd1 _24227_/A sky130_fd_sc_hd__and2_1
X_21438_ _21438_/A vssd1 vssd1 vccd1 vccd1 _21438_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21369_ _21357_/X _21358_/X _21359_/X _21360_/X _21361_/X _21362_/X vssd1 vssd1 vccd1
+ vccd1 _21370_/A sky130_fd_sc_hd__mux4_1
X_24157_ _24157_/A vssd1 vssd1 vccd1 vccd1 _27350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23108_ _23108_/A vssd1 vssd1 vccd1 vccd1 _27097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24088_ _24088_/A vssd1 vssd1 vccd1 vccd1 _27319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15930_ _15930_/A vssd1 vssd1 vccd1 vccd1 _15930_/Y sky130_fd_sc_hd__inv_2
X_27916_ _27916_/A _15988_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
X_23039_ _23107_/S vssd1 vssd1 vccd1 vccd1 _23048_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27847_ _27849_/CLK _27847_/D vssd1 vssd1 vccd1 vccd1 _27847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15861_ _15862_/A vssd1 vssd1 vccd1 vccd1 _15861_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_1103 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _17600_/A vssd1 vssd1 vccd1 vccd1 _25874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14812_ _14812_/A vssd1 vssd1 vccd1 vccd1 _26522_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18580_ _18578_/X _18579_/X _18580_/S vssd1 vssd1 vccd1 vccd1 _18580_/X sky130_fd_sc_hd__mux2_2
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27778_ _27778_/CLK _27778_/D vssd1 vssd1 vccd1 vccd1 _27778_/Q sky130_fd_sc_hd__dfxtp_1
X_15792_ _13072_/X _26102_/Q _15794_/S vssd1 vssd1 vccd1 vccd1 _15793_/A sky130_fd_sc_hd__mux2_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _17599_/S vssd1 vssd1 vccd1 vccd1 _17540_/S sky130_fd_sc_hd__clkbuf_2
X_26729_ _21862_/X _26729_/D vssd1 vssd1 vccd1 vccd1 _26729_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _14743_/A vssd1 vssd1 vccd1 vccd1 _14743_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_550 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17462_ _17462_/A vssd1 vssd1 vccd1 vccd1 _25822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14674_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14686_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16413_ _27384_/Q _16557_/B _16501_/A _14785_/A vssd1 vssd1 vccd1 vccd1 _16413_/X
+ sky130_fd_sc_hd__a22o_1
X_19201_ _19222_/A _19201_/B _19201_/C vssd1 vssd1 vccd1 vccd1 _19202_/A sky130_fd_sc_hd__and3_1
X_13625_ _26924_/Q _13613_/X _13616_/X _13624_/Y vssd1 vssd1 vccd1 vccd1 _26924_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17393_ _20792_/A vssd1 vssd1 vccd1 vccd1 _25655_/A sky130_fd_sc_hd__buf_4
XFILLER_186_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19132_ _26950_/Q _26918_/Q _26886_/Q _26854_/Q _19061_/X _18898_/X vssd1 vssd1 vccd1
+ vccd1 _19132_/X sky130_fd_sc_hd__mux4_2
XFILLER_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16344_ _16242_/S _16182_/X _16185_/X _16186_/X _16369_/A vssd1 vssd1 vccd1 vccd1
+ _16345_/B sky130_fd_sc_hd__o311a_1
X_13556_ _13926_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13556_/Y sky130_fd_sc_hd__nor2_1
Xrepeater76 _27436_/CLK vssd1 vssd1 vccd1 vccd1 _27435_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_158_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater87 _27422_/CLK vssd1 vssd1 vccd1 vccd1 _27293_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater98 _27294_/CLK vssd1 vssd1 vccd1 vccd1 _27121_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_157_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19063_ _27802_/Q _26563_/Q _26435_/Q _26115_/Q _18900_/X _18901_/X vssd1 vssd1 vccd1
+ vccd1 _19063_/X sky130_fd_sc_hd__mux4_2
XFILLER_125_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16275_ _27394_/Q vssd1 vssd1 vccd1 vccd1 _16508_/A sky130_fd_sc_hd__inv_2
XFILLER_160_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ _13558_/A vssd1 vssd1 vccd1 vccd1 _13487_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18014_ _18014_/A vssd1 vssd1 vccd1 vccd1 _18014_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15226_ _14759_/X _26346_/Q _15234_/S vssd1 vssd1 vccd1 vccd1 _15227_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15157_ _15157_/A vssd1 vssd1 vccd1 vccd1 _26377_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _14372_/A _14112_/B vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19965_ _19965_/A vssd1 vssd1 vccd1 vccd1 _19965_/X sky130_fd_sc_hd__clkbuf_1
X_15088_ _14769_/X _26407_/Q _15090_/S vssd1 vssd1 vccd1 vccd1 _15089_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14039_ _14511_/A vssd1 vssd1 vccd1 vccd1 _14399_/A sky130_fd_sc_hd__clkbuf_2
X_18916_ _26813_/Q _26781_/Q _26749_/Q _26717_/Q _18913_/X _24400_/A vssd1 vssd1 vccd1
+ vccd1 _18916_/X sky130_fd_sc_hd__mux4_1
XFILLER_141_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19896_ _19882_/X _19883_/X _19884_/X _19885_/X _19886_/X _19887_/X vssd1 vssd1 vccd1
+ vccd1 _19897_/A sky130_fd_sc_hd__mux4_1
XFILLER_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18847_ _18913_/A vssd1 vssd1 vccd1 vccd1 _18847_/X sky130_fd_sc_hd__buf_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18778_ _18913_/A vssd1 vssd1 vccd1 vccd1 _18778_/X sky130_fd_sc_hd__buf_6
X_17729_ _25928_/Q _17728_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17730_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20740_ _20772_/A vssd1 vssd1 vccd1 vccd1 _20740_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20671_ _20687_/A vssd1 vssd1 vccd1 vccd1 _20671_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22410_ _22410_/A vssd1 vssd1 vccd1 vccd1 _22410_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23390_ _27774_/Q vssd1 vssd1 vccd1 vccd1 _24790_/A sky130_fd_sc_hd__inv_2
XFILLER_148_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22341_ _22331_/X _22332_/X _22333_/X _22334_/X _22335_/X _22336_/X vssd1 vssd1 vccd1
+ vccd1 _22342_/A sky130_fd_sc_hd__mux4_1
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22272_ _22272_/A vssd1 vssd1 vccd1 vccd1 _22272_/X sky130_fd_sc_hd__clkbuf_1
X_25060_ _25060_/A vssd1 vssd1 vccd1 vccd1 _27681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24011_ _24009_/X _24010_/X _24033_/S vssd1 vssd1 vccd1 vccd1 _24011_/X sky130_fd_sc_hd__mux2_1
X_21223_ _21211_/X _21212_/X _21213_/X _21214_/X _21216_/X _21218_/X vssd1 vssd1 vccd1
+ vccd1 _21224_/A sky130_fd_sc_hd__mux4_1
XFILLER_176_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_511 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21154_ _21154_/A vssd1 vssd1 vccd1 vccd1 _21154_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20105_ _20105_/A vssd1 vssd1 vccd1 vccd1 _20105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25962_ _17407_/Y _25962_/D vssd1 vssd1 vccd1 vccd1 _25962_/Q sky130_fd_sc_hd__dfxtp_1
X_21085_ _21077_/X _21078_/X _21079_/X _21080_/X _21081_/X _21082_/X vssd1 vssd1 vccd1
+ vccd1 _21086_/A sky130_fd_sc_hd__mux4_1
XFILLER_144_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27701_ _27703_/CLK _27701_/D vssd1 vssd1 vccd1 vccd1 _27701_/Q sky130_fd_sc_hd__dfxtp_1
X_24913_ _24913_/A _24913_/B vssd1 vssd1 vccd1 vccd1 _24913_/Y sky130_fd_sc_hd__nand2_1
X_20036_ _20028_/X _20029_/X _20030_/X _20031_/X _20032_/X _20033_/X vssd1 vssd1 vccd1
+ vccd1 _20037_/A sky130_fd_sc_hd__mux4_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25893_ _27148_/CLK _25893_/D vssd1 vssd1 vccd1 vccd1 _25893_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27632_ _27633_/CLK _27632_/D vssd1 vssd1 vccd1 vccd1 _27632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24844_ _24844_/A _24844_/B vssd1 vssd1 vccd1 vccd1 _24845_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27563_ _27563_/CLK _27563_/D vssd1 vssd1 vccd1 vccd1 _27563_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24775_ _24803_/A vssd1 vssd1 vccd1 vccd1 _24786_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_21987_ _21981_/X _21982_/X _21983_/X _21984_/X _21985_/X _21986_/X vssd1 vssd1 vccd1
+ vccd1 _21988_/A sky130_fd_sc_hd__mux4_1
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26514_ _21108_/X _26514_/D vssd1 vssd1 vccd1 vccd1 _26514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23726_ _23726_/A vssd1 vssd1 vccd1 vccd1 _27265_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27494_ _27495_/CLK _27494_/D vssd1 vssd1 vccd1 vccd1 _27494_/Q sky130_fd_sc_hd__dfxtp_1
X_20938_ _20954_/A vssd1 vssd1 vccd1 vccd1 _20938_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26445_ _20876_/X _26445_/D vssd1 vssd1 vccd1 vccd1 _26445_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23657_ _24831_/B _27235_/Q _23661_/S vssd1 vssd1 vccd1 vccd1 _23658_/A sky130_fd_sc_hd__mux2_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20869_ _21215_/A vssd1 vssd1 vccd1 vccd1 _20941_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_202_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13410_ _13410_/A vssd1 vssd1 vccd1 vccd1 _26974_/D sky130_fd_sc_hd__clkbuf_1
X_22608_ _22608_/A vssd1 vssd1 vccd1 vccd1 _22608_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14390_ _14390_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _14390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26376_ _20629_/X _26376_/D vssd1 vssd1 vccd1 vccd1 _26376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23588_ _24925_/A _27217_/Q _23595_/S vssd1 vssd1 vccd1 vccd1 _23589_/B sky130_fd_sc_hd__mux2_1
XFILLER_195_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25327_ _27716_/Q _25308_/X _25326_/Y _25297_/X vssd1 vssd1 vccd1 vccd1 _27716_/D
+ sky130_fd_sc_hd__o211a_1
X_13341_ _14731_/A vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__clkbuf_4
X_22539_ _22609_/A vssd1 vssd1 vccd1 vccd1 _22539_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16060_ _27478_/Q _27270_/Q vssd1 vssd1 vccd1 vccd1 _16060_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25258_ _25267_/B _25258_/B vssd1 vssd1 vccd1 vccd1 _25265_/B sky130_fd_sc_hd__or2_1
X_13272_ _27023_/Q _13116_/X _13280_/S vssd1 vssd1 vccd1 vccd1 _13273_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _15749_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _15011_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_679 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24209_ _24209_/A _24210_/B vssd1 vssd1 vccd1 vccd1 _27373_/D sky130_fd_sc_hd__nor2_1
XFILLER_135_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25189_ _25170_/A _25173_/B _25179_/B _25169_/Y vssd1 vssd1 vccd1 vccd1 _25190_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_163_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19750_ _19836_/A vssd1 vssd1 vccd1 vccd1 _19815_/A sky130_fd_sc_hd__clkbuf_2
X_16962_ _27591_/Q vssd1 vssd1 vccd1 vccd1 _16979_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18701_ _18701_/A vssd1 vssd1 vccd1 vccd1 _26013_/D sky130_fd_sc_hd__clkbuf_1
X_15913_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15918_/A sky130_fd_sc_hd__buf_8
X_19681_ _19729_/A vssd1 vssd1 vccd1 vccd1 _19681_/X sky130_fd_sc_hd__clkbuf_1
X_16893_ _16772_/A _16479_/A _16892_/X vssd1 vssd1 vccd1 vccd1 _16893_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18632_ _18689_/S vssd1 vssd1 vccd1 vccd1 _18641_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15844_ _15844_/A vssd1 vssd1 vccd1 vccd1 _26079_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _15775_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15775_/Y sky130_fd_sc_hd__nor2_1
X_18563_ _18557_/X _18559_/X _18562_/X _18150_/A _18489_/X vssd1 vssd1 vccd1 vccd1
+ _18564_/C sky130_fd_sc_hd__a221o_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _27804_/Q _12987_/B vssd1 vssd1 vccd1 vccd1 _12988_/A sky130_fd_sc_hd__and2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17514_ _27436_/Q vssd1 vssd1 vccd1 vccd1 _17514_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14726_/A vssd1 vssd1 vccd1 vccd1 _26549_/D sky130_fd_sc_hd__clkbuf_1
X_18494_ _26965_/Q _26933_/Q _26901_/Q _26869_/Q _18403_/X _18427_/X vssd1 vssd1 vccd1
+ vccd1 _18494_/X sky130_fd_sc_hd__mux4_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _17444_/X _25817_/Q _17454_/S vssd1 vssd1 vccd1 vccd1 _17446_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14657_ _26574_/Q _14645_/X _14653_/X _14656_/Y vssd1 vssd1 vccd1 vccd1 _26574_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13608_ _13878_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13608_/Y sky130_fd_sc_hd__nor2_1
X_17376_ _17374_/X _17375_/X _17386_/S vssd1 vssd1 vccd1 vccd1 _17376_/X sky130_fd_sc_hd__mux2_2
XFILLER_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14588_ _26599_/Q _14576_/X _14579_/X _14587_/Y vssd1 vssd1 vccd1 vccd1 _26599_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19115_ _18996_/X _19114_/X _19089_/X vssd1 vssd1 vccd1 vccd1 _19115_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16327_ _16756_/A vssd1 vssd1 vccd1 vccd1 _16755_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13539_ _26948_/Q _13535_/X _13528_/X _13538_/Y vssd1 vssd1 vccd1 vccd1 _26948_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_199_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19046_ _27801_/Q _26562_/Q _26434_/Q _26114_/Q _18974_/X _19019_/X vssd1 vssd1 vccd1
+ vccd1 _19046_/X sky130_fd_sc_hd__mux4_2
XFILLER_145_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16258_ _27395_/Q vssd1 vssd1 vccd1 vccd1 _16502_/A sky130_fd_sc_hd__inv_2
XFILLER_51_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15209_ _15209_/A vssd1 vssd1 vccd1 vccd1 _26354_/D sky130_fd_sc_hd__clkbuf_1
X_16189_ _27378_/Q vssd1 vssd1 vccd1 vccd1 _23182_/B sky130_fd_sc_hd__inv_2
XFILLER_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28017__483 vssd1 vssd1 vccd1 vccd1 _28017__483/HI _28017_/A sky130_fd_sc_hd__conb_1
X_19948_ _19940_/X _19941_/X _19942_/X _19943_/X _19944_/X _19945_/X vssd1 vssd1 vccd1
+ vccd1 _19949_/A sky130_fd_sc_hd__mux4_1
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19879_ _19879_/A vssd1 vssd1 vccd1 vccd1 _19879_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21910_ _21910_/A vssd1 vssd1 vccd1 vccd1 _21910_/X sky130_fd_sc_hd__clkbuf_1
X_22890_ _22956_/A vssd1 vssd1 vccd1 vccd1 _22890_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21841_ _21825_/X _21826_/X _21827_/X _21828_/X _21830_/X _21832_/X vssd1 vssd1 vccd1
+ vccd1 _21842_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24560_ _24560_/A vssd1 vssd1 vccd1 vccd1 _27541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21772_ _21772_/A vssd1 vssd1 vccd1 vccd1 _21772_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23511_ _23526_/A _23511_/B vssd1 vssd1 vccd1 vccd1 _23512_/A sky130_fd_sc_hd__and2_1
XFILLER_12_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20723_ _20771_/A vssd1 vssd1 vccd1 vccd1 _20723_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24491_ _24635_/B _27581_/Q _27580_/Q _24491_/D vssd1 vssd1 vccd1 vccd1 _24551_/S
+ sky130_fd_sc_hd__and4b_2
XFILLER_51_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26230_ _20121_/X _26230_/D vssd1 vssd1 vccd1 vccd1 _26230_/Q sky130_fd_sc_hd__dfxtp_1
X_23442_ _23482_/A vssd1 vssd1 vccd1 vccd1 _23442_/X sky130_fd_sc_hd__clkbuf_2
X_20654_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20654_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26161_ _19875_/X _26161_/D vssd1 vssd1 vccd1 vccd1 _26161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23373_ _24767_/A _27246_/Q _27253_/Q _24786_/A _23372_/X vssd1 vssd1 vccd1 vccd1
+ _23373_/X sky130_fd_sc_hd__a221o_1
X_20585_ _20601_/A vssd1 vssd1 vccd1 vccd1 _20585_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25112_ _25356_/A vssd1 vssd1 vccd1 vccd1 _25112_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22324_ _22324_/A vssd1 vssd1 vccd1 vccd1 _22324_/X sky130_fd_sc_hd__clkbuf_1
X_26092_ _19632_/X _26092_/D vssd1 vssd1 vccd1 vccd1 _26092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25043_ _25043_/A vssd1 vssd1 vccd1 vccd1 _27679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22255_ _22245_/X _22246_/X _22247_/X _22248_/X _22249_/X _22250_/X vssd1 vssd1 vccd1
+ vccd1 _22256_/A sky130_fd_sc_hd__mux4_1
XFILLER_180_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21206_ _21206_/A vssd1 vssd1 vccd1 vccd1 _21206_/X sky130_fd_sc_hd__clkbuf_1
X_22186_ _22186_/A vssd1 vssd1 vccd1 vccd1 _22186_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21137_ _21125_/X _21126_/X _21127_/X _21128_/X _21130_/X _21132_/X vssd1 vssd1 vccd1
+ vccd1 _21138_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26994_ _22782_/X _26994_/D vssd1 vssd1 vccd1 vccd1 _26994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21068_ _21068_/A vssd1 vssd1 vccd1 vccd1 _21068_/X sky130_fd_sc_hd__clkbuf_1
X_25945_ _27312_/CLK _25945_/D vssd1 vssd1 vccd1 vccd1 _25945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20019_ _20019_/A vssd1 vssd1 vccd1 vccd1 _20019_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _26830_/Q _13880_/X _13886_/X _13889_/Y vssd1 vssd1 vccd1 vccd1 _26830_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25876_ _27827_/CLK _25876_/D vssd1 vssd1 vccd1 vccd1 _25876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27615_ _27617_/CLK _27615_/D vssd1 vssd1 vccd1 vccd1 _27615_/Q sky130_fd_sc_hd__dfxtp_1
X_24827_ _27642_/Q _25564_/A _24733_/Y vssd1 vssd1 vccd1 vccd1 _24828_/C sky130_fd_sc_hd__a21bo_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27546_ _27568_/CLK _27546_/D vssd1 vssd1 vccd1 vccd1 _27546_/Q sky130_fd_sc_hd__dfxtp_1
X_15560_ _26198_/Q _14721_/A _15562_/S vssd1 vssd1 vccd1 vccd1 _15561_/A sky130_fd_sc_hd__mux2_1
X_24758_ _24771_/A vssd1 vssd1 vccd1 vccd1 _24758_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14511_ _14511_/A vssd1 vssd1 vccd1 vccd1 _15767_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23709_ _23709_/A vssd1 vssd1 vccd1 vccd1 _27258_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27477_ _27477_/CLK _27477_/D vssd1 vssd1 vccd1 vccd1 _27477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15491_ _15491_/A vssd1 vssd1 vccd1 vccd1 _26229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24689_ _27177_/Q _24698_/B vssd1 vssd1 vccd1 vccd1 _24689_/X sky130_fd_sc_hd__or2_1
XFILLER_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17230_ _17291_/A vssd1 vssd1 vccd1 vccd1 _17280_/S sky130_fd_sc_hd__buf_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14442_ _16298_/A vssd1 vssd1 vccd1 vccd1 _15716_/A sky130_fd_sc_hd__buf_2
X_26428_ _20813_/X _26428_/D vssd1 vssd1 vccd1 vccd1 _26428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17161_ _17116_/X _17154_/X _17157_/X _17160_/X vssd1 vssd1 vccd1 vccd1 _17161_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_196_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14373_ _26666_/Q _14365_/X _14371_/X _14372_/Y vssd1 vssd1 vccd1 vccd1 _26666_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26359_ _20565_/X _26359_/D vssd1 vssd1 vccd1 vccd1 _26359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16112_ _16112_/A _16112_/B vssd1 vssd1 vccd1 vccd1 _16201_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ _13324_/A vssd1 vssd1 vccd1 vccd1 _27001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17092_ _17092_/A vssd1 vssd1 vccd1 vccd1 _27922_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16043_ _27476_/Q _27372_/Q vssd1 vssd1 vccd1 vccd1 _16043_/Y sky130_fd_sc_hd__nand2_1
X_13255_ _13255_/A vssd1 vssd1 vccd1 vccd1 _27031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _13186_/A vssd1 vssd1 vccd1 vccd1 _27043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19802_ _19796_/X _19797_/X _19798_/X _19799_/X _19800_/X _19801_/X vssd1 vssd1 vccd1
+ vccd1 _19803_/A sky130_fd_sc_hd__mux4_1
XFILLER_111_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17994_ _18443_/A vssd1 vssd1 vccd1 vccd1 _18468_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19733_ _19801_/A vssd1 vssd1 vccd1 vccd1 _19733_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16945_ _16945_/A _16945_/B _16945_/C vssd1 vssd1 vccd1 vccd1 _16945_/X sky130_fd_sc_hd__and3_1
XFILLER_77_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19664_ _19836_/A vssd1 vssd1 vccd1 vccd1 _19729_/A sky130_fd_sc_hd__clkbuf_2
X_16876_ _24253_/A _24245_/A _24243_/A _16875_/X vssd1 vssd1 vccd1 vccd1 _16896_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18615_ _27690_/Q _18591_/X _18594_/X _18614_/Y vssd1 vssd1 vccd1 vccd1 _18615_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _13166_/X _26086_/Q _15827_/S vssd1 vssd1 vccd1 vccd1 _15828_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19595_ _19589_/X _19590_/X _19591_/X _19592_/X _19593_/X _19594_/X vssd1 vssd1 vccd1
+ vccd1 _19596_/A sky130_fd_sc_hd__mux4_1
X_15758_ _15758_/A _15758_/B vssd1 vssd1 vccd1 vccd1 _15758_/Y sky130_fd_sc_hd__nor2_1
X_18546_ _18842_/A _18546_/B _18546_/C vssd1 vssd1 vccd1 vccd1 _18547_/A sky130_fd_sc_hd__and3_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14709_ _14709_/A vssd1 vssd1 vccd1 vccd1 _14709_/X sky130_fd_sc_hd__buf_2
X_18477_ _18468_/X _18471_/X _18476_/X _18412_/X vssd1 vssd1 vccd1 vccd1 _18491_/B
+ sky130_fd_sc_hd__a211o_1
X_15689_ _13228_/X _26140_/Q _15689_/S vssd1 vssd1 vccd1 vccd1 _15690_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17428_ _27409_/Q vssd1 vssd1 vccd1 vccd1 _17428_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ _27855_/Q _27159_/Q _25904_/Q _25872_/Q _17325_/X _17313_/X vssd1 vssd1 vccd1
+ vccd1 _17359_/X sky130_fd_sc_hd__mux4_1
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20370_ _20354_/X _20357_/X _20360_/X _20363_/X _20364_/X _20365_/X vssd1 vssd1 vccd1
+ vccd1 _20371_/A sky130_fd_sc_hd__mux4_1
XFILLER_174_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19029_ _26273_/Q _26241_/Q _26209_/Q _26177_/Q _19028_/X _18955_/X vssd1 vssd1 vccd1
+ vccd1 _19029_/X sky130_fd_sc_hd__mux4_2
XFILLER_106_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22040_ _22072_/A vssd1 vssd1 vccd1 vccd1 _22040_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23991_ _23991_/A vssd1 vssd1 vccd1 vccd1 _23991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25730_ _25730_/A vssd1 vssd1 vccd1 vccd1 _25730_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22942_ _22958_/A vssd1 vssd1 vccd1 vccd1 _22942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25661_ _25709_/A vssd1 vssd1 vccd1 vccd1 _25661_/X sky130_fd_sc_hd__clkbuf_2
X_22873_ _22959_/A vssd1 vssd1 vccd1 vccd1 _22943_/A sky130_fd_sc_hd__buf_2
X_27400_ _27404_/CLK _27400_/D vssd1 vssd1 vccd1 vccd1 _27400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24612_ _27665_/Q _24620_/B vssd1 vssd1 vccd1 vccd1 _24613_/A sky130_fd_sc_hd__and2_1
X_21824_ _21824_/A vssd1 vssd1 vccd1 vccd1 _21824_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25592_ _25592_/A vssd1 vssd1 vccd1 vccd1 _25592_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27331_ _27331_/CLK _27331_/D vssd1 vssd1 vccd1 vccd1 _27331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24543_ _24552_/A _24543_/B vssd1 vssd1 vccd1 vccd1 _24544_/A sky130_fd_sc_hd__and2_1
X_21755_ _21737_/X _21738_/X _21739_/X _21740_/X _21743_/X _21746_/X vssd1 vssd1 vccd1
+ vccd1 _21756_/A sky130_fd_sc_hd__mux4_1
XFILLER_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20706_ _20706_/A vssd1 vssd1 vccd1 vccd1 _20772_/A sky130_fd_sc_hd__buf_2
X_27262_ _27262_/CLK _27262_/D vssd1 vssd1 vccd1 vccd1 _27262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24474_ _27634_/Q _24478_/B vssd1 vssd1 vccd1 vccd1 _24475_/A sky130_fd_sc_hd__and2_1
XFILLER_197_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21686_ _21686_/A vssd1 vssd1 vccd1 vccd1 _21686_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26213_ _20057_/X _26213_/D vssd1 vssd1 vccd1 vccd1 _26213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23425_ _27164_/Q _23430_/B vssd1 vssd1 vccd1 vccd1 _23425_/X sky130_fd_sc_hd__or2_1
X_27193_ _27536_/CLK _27193_/D vssd1 vssd1 vccd1 vccd1 _27193_/Q sky130_fd_sc_hd__dfxtp_1
X_20637_ _20685_/A vssd1 vssd1 vccd1 vccd1 _20637_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26144_ _19811_/X _26144_/D vssd1 vssd1 vccd1 vccd1 _26144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23356_ _27763_/Q vssd1 vssd1 vccd1 vccd1 _24759_/A sky130_fd_sc_hd__clkinv_2
X_20568_ _20600_/A vssd1 vssd1 vccd1 vccd1 _20568_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22307_ _22299_/X _22300_/X _22301_/X _22302_/X _22303_/X _22304_/X vssd1 vssd1 vccd1
+ vccd1 _22308_/A sky130_fd_sc_hd__mux4_1
XFILLER_109_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26075_ _19580_/X _26075_/D vssd1 vssd1 vccd1 vccd1 _26075_/Q sky130_fd_sc_hd__dfxtp_1
X_23287_ _27732_/Q _23284_/Y _27744_/Q _23285_/Y _23286_/X vssd1 vssd1 vccd1 vccd1
+ _23293_/B sky130_fd_sc_hd__a221o_1
XFILLER_164_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20499_ _20515_/A vssd1 vssd1 vccd1 vccd1 _20499_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ _16017_/B vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__clkbuf_2
X_25026_ _27832_/Q _27136_/Q _25881_/Q _25849_/Q _25018_/X _24991_/X vssd1 vssd1 vccd1
+ vccd1 _25026_/X sky130_fd_sc_hd__mux4_1
X_22238_ _22238_/A vssd1 vssd1 vccd1 vccd1 _22238_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22169_ _22157_/X _22158_/X _22159_/X _22160_/X _22161_/X _22162_/X vssd1 vssd1 vccd1
+ vccd1 _22170_/A sky130_fd_sc_hd__mux4_1
XFILLER_160_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14991_ _26447_/Q _14988_/X _14989_/X _14990_/Y vssd1 vssd1 vccd1 vccd1 _26447_/D
+ sky130_fd_sc_hd__a31o_1
X_26977_ _22730_/X _26977_/D vssd1 vssd1 vccd1 vccd1 _26977_/Q sky130_fd_sc_hd__dfxtp_1
X_13942_ _14813_/B _14149_/B vssd1 vssd1 vccd1 vccd1 _13964_/A sky130_fd_sc_hd__or2_1
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16730_ _16726_/Y _16727_/X _16728_/X _16729_/X vssd1 vssd1 vccd1 vccd1 _24233_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_25928_ _27844_/CLK _25928_/D vssd1 vssd1 vccd1 vccd1 _25928_/Q sky130_fd_sc_hd__dfxtp_1
X_16661_ _16660_/Y _16885_/B _16548_/Y vssd1 vssd1 vccd1 vccd1 _16662_/B sky130_fd_sc_hd__o21bai_1
X_13873_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13873_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25859_ _27844_/CLK _25859_/D vssd1 vssd1 vccd1 vccd1 _25859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15612_ _15612_/A vssd1 vssd1 vccd1 vccd1 _26175_/D sky130_fd_sc_hd__clkbuf_1
X_18400_ _18844_/A vssd1 vssd1 vccd1 vccd1 _18509_/A sky130_fd_sc_hd__clkbuf_1
X_16592_ _16791_/B vssd1 vssd1 vccd1 vccd1 _16599_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19380_ _18801_/X _19375_/X _19377_/X _19379_/X _19360_/X vssd1 vssd1 vccd1 vccd1
+ _19381_/C sky130_fd_sc_hd__a221o_1
XFILLER_131_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _18328_/X _18330_/X _18331_/S vssd1 vssd1 vccd1 vccd1 _18331_/X sky130_fd_sc_hd__mux2_2
X_15543_ _13222_/X _26205_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15544_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27529_ _27529_/CLK _27529_/D vssd1 vssd1 vccd1 vccd1 _27529_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18260_/X _18261_/X _18331_/S vssd1 vssd1 vccd1 vccd1 _18262_/X sky130_fd_sc_hd__mux2_1
X_15474_ _15474_/A vssd1 vssd1 vccd1 vccd1 _26236_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17213_ _27211_/Q _17212_/X _17250_/S vssd1 vssd1 vccd1 vccd1 _17214_/A sky130_fd_sc_hd__mux2_1
X_14425_ _14425_/A vssd1 vssd1 vccd1 vccd1 _15703_/A sky130_fd_sc_hd__buf_2
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18193_ _18264_/A _18193_/B _18193_/C vssd1 vssd1 vccd1 vccd1 _18194_/A sky130_fd_sc_hd__and3_1
XFILLER_168_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17144_ _17266_/A vssd1 vssd1 vccd1 vccd1 _17193_/S sky130_fd_sc_hd__clkbuf_2
X_14356_ _14356_/A _14363_/B vssd1 vssd1 vccd1 vccd1 _14356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ _27007_/Q _13210_/X _13313_/S vssd1 vssd1 vccd1 vccd1 _13308_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17075_ _17052_/X _17070_/X _17072_/X _17074_/X vssd1 vssd1 vccd1 vccd1 _17075_/X
+ sky130_fd_sc_hd__o22a_1
X_14287_ _14374_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16026_ _16297_/B _16296_/B _26073_/Q vssd1 vssd1 vccd1 vccd1 _16026_/X sky130_fd_sc_hd__or3b_1
XFILLER_157_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13238_ _27335_/Q _13193_/X _13194_/X _27303_/Q _13237_/X vssd1 vssd1 vccd1 vccd1
+ _16182_/A sky130_fd_sc_hd__a221o_1
XFILLER_143_469 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13169_ _27282_/Q _13169_/B vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__and2_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17977_ _26687_/Q _26655_/Q _26623_/Q _26591_/Q _17865_/X _17928_/X vssd1 vssd1 vccd1
+ vccd1 _17979_/A sky130_fd_sc_hd__mux4_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19716_ _19710_/X _19711_/X _19712_/X _19713_/X _19714_/X _19715_/X vssd1 vssd1 vccd1
+ vccd1 _19717_/A sky130_fd_sc_hd__mux4_1
X_16928_ _27486_/Q vssd1 vssd1 vccd1 vccd1 _24208_/A sky130_fd_sc_hd__inv_2
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19647_ _19715_/A vssd1 vssd1 vccd1 vccd1 _19647_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16859_ _25909_/Q _16752_/A _16754_/A _16646_/B vssd1 vssd1 vccd1 vccd1 _16859_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19578_ _19626_/A vssd1 vssd1 vccd1 vccd1 _19578_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18529_ _18529_/A vssd1 vssd1 vccd1 vccd1 _25972_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21540_ _21540_/A vssd1 vssd1 vccd1 vccd1 _21540_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21471_ _21459_/X _21460_/X _21461_/X _21462_/X _21463_/X _21464_/X vssd1 vssd1 vccd1
+ vccd1 _21472_/A sky130_fd_sc_hd__mux4_1
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23210_ _23210_/A vssd1 vssd1 vccd1 vccd1 _27141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20422_ _20408_/X _20409_/X _20410_/X _20411_/X _20412_/X _20413_/X vssd1 vssd1 vccd1
+ vccd1 _20423_/A sky130_fd_sc_hd__mux4_1
XFILLER_181_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24190_ _24190_/A vssd1 vssd1 vccd1 vccd1 _27365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23141_ _27111_/Q _17718_/X _23143_/S vssd1 vssd1 vccd1 vccd1 _23142_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20353_ _20702_/A vssd1 vssd1 vccd1 vccd1 _20424_/A sky130_fd_sc_hd__buf_2
XFILLER_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23072_ _23094_/A vssd1 vssd1 vccd1 vccd1 _23081_/S sky130_fd_sc_hd__clkbuf_2
X_20284_ _20267_/X _20269_/X _20271_/X _20273_/X _20274_/X _20275_/X vssd1 vssd1 vccd1
+ vccd1 _20285_/A sky130_fd_sc_hd__mux4_1
XFILLER_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22023_ _22071_/A vssd1 vssd1 vccd1 vccd1 _22023_/X sky130_fd_sc_hd__clkbuf_2
X_26900_ _22462_/X _26900_/D vssd1 vssd1 vccd1 vccd1 _26900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26831_ _22222_/X _26831_/D vssd1 vssd1 vccd1 vccd1 _26831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26762_ _21976_/X _26762_/D vssd1 vssd1 vccd1 vccd1 _26762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23974_ _23943_/X _23972_/X _23973_/X _23958_/X vssd1 vssd1 vccd1 vccd1 _27293_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25713_ _25705_/X _25706_/X _25707_/X _25708_/X _25709_/X _25710_/X vssd1 vssd1 vccd1
+ vccd1 _25714_/A sky130_fd_sc_hd__mux4_1
X_22925_ _22957_/A vssd1 vssd1 vccd1 vccd1 _22925_/X sky130_fd_sc_hd__clkbuf_1
X_26693_ _21734_/X _26693_/D vssd1 vssd1 vccd1 vccd1 _26693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25644_ _25644_/A vssd1 vssd1 vccd1 vccd1 _25644_/X sky130_fd_sc_hd__clkbuf_1
X_22856_ _22872_/A vssd1 vssd1 vccd1 vccd1 _22856_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21807_ _21793_/X _21794_/X _21795_/X _21796_/X _21797_/X _21798_/X vssd1 vssd1 vccd1
+ vccd1 _21808_/A sky130_fd_sc_hd__mux4_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25575_ _27712_/Q _25568_/X _25569_/X vssd1 vssd1 vccd1 vccd1 _25575_/Y sky130_fd_sc_hd__a21oi_1
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22787_ _22959_/A vssd1 vssd1 vccd1 vccd1 _22857_/A sky130_fd_sc_hd__clkbuf_2
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27314_ _27388_/CLK _27314_/D vssd1 vssd1 vccd1 vccd1 _27314_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24526_ _24524_/X _24525_/X _24499_/X vssd1 vssd1 vccd1 vccd1 _27530_/D sky130_fd_sc_hd__o21a_1
X_21738_ _21738_/A vssd1 vssd1 vccd1 vccd1 _21738_/X sky130_fd_sc_hd__clkbuf_1
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27245_ _27245_/CLK _27245_/D vssd1 vssd1 vccd1 vccd1 _27245_/Q sky130_fd_sc_hd__dfxtp_1
X_24457_ _24457_/A vssd1 vssd1 vccd1 vccd1 _27505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21669_ _22017_/A vssd1 vssd1 vccd1 vccd1 _21738_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14210_ _14388_/A _14213_/B vssd1 vssd1 vccd1 vccd1 _14210_/Y sky130_fd_sc_hd__nor2_1
X_23408_ _24848_/A _23405_/Y _27247_/Q _24769_/A _23407_/X vssd1 vssd1 vccd1 vccd1
+ _23408_/X sky130_fd_sc_hd__o221a_1
XFILLER_71_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27176_ _27607_/CLK _27176_/D vssd1 vssd1 vccd1 vccd1 _27176_/Q sky130_fd_sc_hd__dfxtp_1
X_15190_ _15190_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15247_/A sky130_fd_sc_hd__or2_4
X_24388_ _24388_/A _24638_/A vssd1 vssd1 vccd1 vccd1 _24389_/A sky130_fd_sc_hd__and2_1
XFILLER_165_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14141_ _26749_/Q _14130_/X _14133_/X _14140_/Y vssd1 vssd1 vccd1 vccd1 _26749_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_153_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26127_ _19759_/X _26127_/D vssd1 vssd1 vccd1 vccd1 _26127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23339_ _24825_/A _27234_/Q _27257_/Q _24796_/A vssd1 vssd1 vccd1 vccd1 _23361_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14072_ _14079_/A vssd1 vssd1 vccd1 vccd1 _14127_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26058_ _26068_/CLK _26058_/D vssd1 vssd1 vccd1 vccd1 _26058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25009_ _27229_/Q vssd1 vssd1 vccd1 vccd1 _25009_/X sky130_fd_sc_hd__buf_2
X_17900_ _17900_/A vssd1 vssd1 vccd1 vccd1 _18486_/A sky130_fd_sc_hd__clkbuf_4
X_13023_ _27368_/Q _27367_/Q vssd1 vssd1 vccd1 vccd1 _13194_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18880_ _19393_/A vssd1 vssd1 vccd1 vccd1 _18880_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17831_ _18360_/A vssd1 vssd1 vccd1 vccd1 _18358_/A sky130_fd_sc_hd__buf_4
XFILLER_126_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17762_ _17762_/A vssd1 vssd1 vccd1 vccd1 _25938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14974_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19501_ _19501_/A _19501_/B vssd1 vssd1 vccd1 vccd1 _19501_/X sky130_fd_sc_hd__or2_1
XFILLER_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16713_ _16774_/A _16711_/Y _16712_/X vssd1 vssd1 vccd1 vccd1 _16713_/Y sky130_fd_sc_hd__o21ai_1
X_13925_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13925_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17693_ _17776_/S vssd1 vssd1 vccd1 vccd1 _17706_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_48_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19432_ _26707_/Q _26675_/Q _26643_/Q _26611_/Q _19317_/X _19385_/X vssd1 vssd1 vccd1
+ vccd1 _19432_/X sky130_fd_sc_hd__mux4_2
X_13856_ _13872_/A vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16644_ _16583_/A _16831_/B _16643_/X vssd1 vssd1 vccd1 vccd1 _16644_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19363_ _19363_/A vssd1 vssd1 vccd1 vccd1 _26063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13787_ _13827_/A vssd1 vssd1 vccd1 vccd1 _13799_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16575_ _25971_/Q _16098_/X _16574_/X vssd1 vssd1 vccd1 vccd1 _16916_/A sky130_fd_sc_hd__a21oi_4
XFILLER_188_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18314_ _18312_/X _18313_/X _18378_/S vssd1 vssd1 vccd1 vccd1 _18314_/X sky130_fd_sc_hd__mux2_1
X_15526_ _13172_/X _26213_/Q _15534_/S vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__mux2_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _26957_/Q _26925_/Q _26893_/Q _26861_/Q _18913_/A _19445_/A vssd1 vssd1 vccd1
+ vccd1 _19294_/X sky130_fd_sc_hd__mux4_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18245_ _26954_/Q _26922_/Q _26890_/Q _26858_/Q _18244_/X _18129_/X vssd1 vssd1 vccd1
+ vccd1 _18245_/X sky130_fd_sc_hd__mux4_2
X_15457_ _15457_/A vssd1 vssd1 vccd1 vccd1 _26244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14408_ _14408_/A _14412_/B vssd1 vssd1 vccd1 vccd1 _14408_/Y sky130_fd_sc_hd__nor2_1
XFILLER_198_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18176_ _26823_/Q _26791_/Q _26759_/Q _26727_/Q _18175_/X _18058_/X vssd1 vssd1 vccd1
+ vccd1 _18176_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15388_ _14785_/X _26274_/Q _15390_/S vssd1 vssd1 vccd1 vccd1 _15389_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ _14393_/A vssd1 vssd1 vccd1 vccd1 _14350_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17127_ _17123_/X _17125_/X _17174_/S vssd1 vssd1 vccd1 vccd1 _17127_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17058_ _25815_/Q _26014_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17058_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16009_ _16132_/A vssd1 vssd1 vccd1 vccd1 _16264_/B sky130_fd_sc_hd__clkbuf_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater300 _27654_/CLK vssd1 vssd1 vccd1 vccd1 _27658_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater311 _27542_/CLK vssd1 vssd1 vccd1 vccd1 _27472_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater322 _27711_/CLK vssd1 vssd1 vccd1 vccd1 _27629_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater333 _27772_/CLK vssd1 vssd1 vccd1 vccd1 _27768_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater344 _27642_/CLK vssd1 vssd1 vccd1 vccd1 _27690_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater355 _27575_/CLK vssd1 vssd1 vccd1 vccd1 _27569_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater366 _27411_/CLK vssd1 vssd1 vccd1 vccd1 _27410_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater377 _27452_/CLK vssd1 vssd1 vccd1 vccd1 _27651_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20971_ _21143_/A vssd1 vssd1 vccd1 vccd1 _21039_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater388 _27196_/CLK vssd1 vssd1 vccd1 vccd1 _27208_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater399 _27576_/CLK vssd1 vssd1 vccd1 vccd1 _27442_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22710_ _22710_/A vssd1 vssd1 vccd1 vccd1 _22710_/X sky130_fd_sc_hd__clkbuf_1
X_23690_ _27770_/Q _27250_/Q _23694_/S vssd1 vssd1 vccd1 vccd1 _23691_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22641_ _22630_/X _22632_/X _22634_/X _22636_/X _22637_/X _22638_/X vssd1 vssd1 vccd1
+ vccd1 _22642_/A sky130_fd_sc_hd__mux4_1
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25360_ _25428_/S vssd1 vssd1 vccd1 vccd1 _25369_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22572_ _22572_/A vssd1 vssd1 vccd1 vccd1 _22572_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24311_ _27540_/Q _24317_/B vssd1 vssd1 vccd1 vccd1 _24312_/A sky130_fd_sc_hd__and2_1
X_21523_ _21513_/X _21514_/X _21515_/X _21516_/X _21517_/X _21518_/X vssd1 vssd1 vccd1
+ vccd1 _21524_/A sky130_fd_sc_hd__mux4_1
XFILLER_194_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25291_ _25306_/A _25291_/B vssd1 vssd1 vccd1 vccd1 _25291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27030_ _22914_/X _27030_/D vssd1 vssd1 vccd1 vccd1 _27030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24242_ _24242_/A _24256_/B vssd1 vssd1 vccd1 vccd1 _27392_/D sky130_fd_sc_hd__nor2_1
X_21454_ _21454_/A vssd1 vssd1 vccd1 vccd1 _21454_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20405_ _20405_/A vssd1 vssd1 vccd1 vccd1 _20405_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24173_ _27463_/Q _24173_/B vssd1 vssd1 vccd1 vccd1 _24174_/A sky130_fd_sc_hd__and2_1
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21385_ _21373_/X _21374_/X _21375_/X _21376_/X _21377_/X _21378_/X vssd1 vssd1 vccd1
+ vccd1 _21386_/A sky130_fd_sc_hd__mux4_1
XFILLER_179_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23124_ _27103_/Q _17692_/X _23132_/S vssd1 vssd1 vccd1 vccd1 _23125_/A sky130_fd_sc_hd__mux2_1
X_20336_ _20336_/A vssd1 vssd1 vccd1 vccd1 _20336_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_406 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27932_ _27932_/A _15953_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23055_ _27073_/Q _17699_/X _23059_/S vssd1 vssd1 vccd1 vccd1 _23056_/A sky130_fd_sc_hd__mux2_1
X_20267_ _20334_/A vssd1 vssd1 vccd1 vccd1 _20267_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22006_ _22006_/A vssd1 vssd1 vccd1 vccd1 _22006_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20198_ _20181_/X _20183_/X _20185_/X _20187_/X _20188_/X _20189_/X vssd1 vssd1 vccd1
+ vccd1 _20199_/A sky130_fd_sc_hd__mux4_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26814_ _22156_/X _26814_/D vssd1 vssd1 vccd1 vccd1 _26814_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27794_ _25630_/X _27794_/D vssd1 vssd1 vccd1 vccd1 _27794_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26745_ _21920_/X _26745_/D vssd1 vssd1 vccd1 vccd1 _26745_/Q sky130_fd_sc_hd__dfxtp_1
X_23957_ _27086_/Q _23954_/X _23955_/X _27118_/Q _23956_/X vssd1 vssd1 vccd1 vccd1
+ _23957_/X sky130_fd_sc_hd__a221o_1
XFILLER_99_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13710_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22908_ _22956_/A vssd1 vssd1 vccd1 vccd1 _22908_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26676_ _21682_/X _26676_/D vssd1 vssd1 vccd1 vccd1 _26676_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _26562_/Q _14685_/X _14679_/X _14689_/Y vssd1 vssd1 vccd1 vccd1 _26562_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23888_ _23849_/X _23886_/X _23887_/X _23864_/X vssd1 vssd1 vccd1 vccd1 _27284_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _26918_/Q _13639_/X _13629_/X _13640_/Y vssd1 vssd1 vccd1 vccd1 _26918_/D
+ sky130_fd_sc_hd__a31o_1
X_22839_ _22871_/A vssd1 vssd1 vccd1 vccd1 _22839_/X sky130_fd_sc_hd__clkbuf_1
X_25627_ _23025_/X _23026_/X _23027_/X _23028_/X _23029_/X _23030_/X vssd1 vssd1 vccd1
+ vccd1 _25628_/A sky130_fd_sc_hd__mux4_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16360_/A _16447_/B vssd1 vssd1 vccd1 vccd1 _16361_/B sky130_fd_sc_hd__nand2_1
X_13572_ _14524_/A vssd1 vssd1 vccd1 vccd1 _13936_/A sky130_fd_sc_hd__clkbuf_2
X_25558_ _24786_/A _25534_/X _25551_/Y _25556_/X _25557_/X vssd1 vssd1 vccd1 vccd1
+ _27773_/D sky130_fd_sc_hd__a221oi_1
XFILLER_13_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15311_ _26308_/Q _13389_/X _15317_/S vssd1 vssd1 vccd1 vccd1 _15312_/A sky130_fd_sc_hd__mux2_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24509_ _27604_/Q _24509_/B vssd1 vssd1 vccd1 vccd1 _24510_/A sky130_fd_sc_hd__and2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16291_ _16802_/A _16623_/B vssd1 vssd1 vccd1 vccd1 _16292_/D sky130_fd_sc_hd__or2b_1
X_25489_ _25470_/X _25182_/B _25488_/X _25483_/X vssd1 vssd1 vccd1 vccd1 _25489_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _15242_/A vssd1 vssd1 vccd1 vccd1 _26339_/D sky130_fd_sc_hd__clkbuf_1
X_18030_ _24611_/A vssd1 vssd1 vccd1 vccd1 _18146_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_157_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27228_ _27790_/CLK _27228_/D vssd1 vssd1 vccd1 vccd1 _27228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27159_ _27855_/CLK _27159_/D vssd1 vssd1 vccd1 vccd1 _27159_/Q sky130_fd_sc_hd__dfxtp_1
X_15173_ _26369_/Q _13398_/X _15173_/S vssd1 vssd1 vccd1 vccd1 _15174_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14124_ _26756_/Q _14117_/X _14120_/X _14123_/Y vssd1 vssd1 vccd1 vccd1 _26756_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_193_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19981_ _19981_/A vssd1 vssd1 vccd1 vccd1 _19981_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ _14527_/A vssd1 vssd1 vccd1 vccd1 _14410_/A sky130_fd_sc_hd__clkbuf_2
X_18932_ _18932_/A vssd1 vssd1 vccd1 vccd1 _18932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ _13006_/A vssd1 vssd1 vccd1 vccd1 _27796_/D sky130_fd_sc_hd__clkbuf_1
X_18863_ _19287_/A vssd1 vssd1 vccd1 vccd1 _18863_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17814_ _17814_/A _17813_/X vssd1 vssd1 vccd1 vccd1 _17814_/X sky130_fd_sc_hd__or2b_1
XFILLER_95_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18794_ _18897_/A vssd1 vssd1 vccd1 vccd1 _19321_/A sky130_fd_sc_hd__buf_2
XFILLER_48_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17745_ _25933_/Q _17744_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17746_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14957_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14957_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _13908_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _13908_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17676_ _17757_/A vssd1 vssd1 vccd1 vccd1 _17776_/S sky130_fd_sc_hd__buf_2
XFILLER_39_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14888_ _14709_/X _26489_/Q _14896_/S vssd1 vssd1 vccd1 vccd1 _14889_/A sky130_fd_sc_hd__mux2_1
X_19415_ _27817_/Q _26578_/Q _26450_/Q _26130_/Q _19414_/X _19321_/X vssd1 vssd1 vccd1
+ vccd1 _19415_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16627_ _16618_/Y _16620_/X _16624_/X _16626_/X vssd1 vssd1 vccd1 vccd1 _24250_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13839_ _26846_/Q _13832_/X _13833_/X _13838_/Y vssd1 vssd1 vccd1 vccd1 _26846_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ _19344_/X _19345_/X _19346_/S vssd1 vssd1 vccd1 vccd1 _19346_/X sky130_fd_sc_hd__mux2_1
X_16558_ _16298_/A _16400_/A _16067_/X _16556_/Y _16557_/Y vssd1 vssd1 vccd1 vccd1
+ _16648_/C sky130_fd_sc_hd__o221a_2
XFILLER_188_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15509_ _15509_/A vssd1 vssd1 vccd1 vccd1 _26221_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19277_ _27811_/Q _26572_/Q _26444_/Q _26124_/Q _19255_/X _19183_/X vssd1 vssd1 vccd1
+ vccd1 _19277_/X sky130_fd_sc_hd__mux4_2
XFILLER_202_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16489_ _16670_/A _16497_/B _16489_/C vssd1 vssd1 vccd1 vccd1 _16493_/C sky130_fd_sc_hd__nand3_1
XFILLER_31_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18228_ _18387_/A vssd1 vssd1 vccd1 vccd1 _18228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _18150_/X _18153_/X _18158_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _18170_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_190_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21170_ _21170_/A vssd1 vssd1 vccd1 vccd1 _21170_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20121_ _20121_/A vssd1 vssd1 vccd1 vccd1 _20121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20052_ _20044_/X _20045_/X _20046_/X _20047_/X _20048_/X _20049_/X vssd1 vssd1 vccd1
+ vccd1 _20053_/A sky130_fd_sc_hd__mux4_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24860_ _27648_/Q _24834_/X _24859_/Y _24839_/X vssd1 vssd1 vccd1 vccd1 _27648_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater130 _26039_/CLK vssd1 vssd1 vccd1 vccd1 _27125_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater141 _27115_/CLK vssd1 vssd1 vccd1 vccd1 _27083_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23811_ _23807_/X _23809_/X _23846_/S vssd1 vssd1 vccd1 vccd1 _23811_/X sky130_fd_sc_hd__mux2_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater152 _27418_/CLK vssd1 vssd1 vccd1 vccd1 _27788_/CLK sky130_fd_sc_hd__clkbuf_1
X_24791_ _27629_/Q _24785_/X _24790_/Y _24787_/X vssd1 vssd1 vccd1 vccd1 _27629_/D
+ sky130_fd_sc_hd__o211a_1
Xrepeater163 _27827_/CLK vssd1 vssd1 vccd1 vccd1 _27132_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater174 _26022_/CLK vssd1 vssd1 vccd1 vccd1 _25925_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater185 _27414_/CLK vssd1 vssd1 vccd1 vccd1 _25917_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26530_ _21170_/X _26530_/D vssd1 vssd1 vccd1 vccd1 _26530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _14507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23742_ _23777_/A vssd1 vssd1 vccd1 vccd1 _23997_/A sky130_fd_sc_hd__buf_2
XFILLER_66_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater196 _27676_/CLK vssd1 vssd1 vccd1 vccd1 _25980_/CLK sky130_fd_sc_hd__clkbuf_1
X_20954_ _20954_/A vssd1 vssd1 vccd1 vccd1 _20954_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_219 _14753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26461_ _20930_/X _26461_/D vssd1 vssd1 vccd1 vccd1 _26461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23673_ _23673_/A vssd1 vssd1 vccd1 vccd1 _27242_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _21143_/A vssd1 vssd1 vccd1 vccd1 _20953_/A sky130_fd_sc_hd__clkbuf_4
X_25412_ _25412_/A vssd1 vssd1 vccd1 vccd1 _27744_/D sky130_fd_sc_hd__clkbuf_1
X_22624_ _22624_/A vssd1 vssd1 vccd1 vccd1 _22624_/X sky130_fd_sc_hd__clkbuf_1
X_26392_ _20679_/X _26392_/D vssd1 vssd1 vccd1 vccd1 _26392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25343_ _25343_/A _25343_/B vssd1 vssd1 vccd1 vccd1 _25344_/B sky130_fd_sc_hd__xor2_2
X_22555_ _22539_/X _22542_/X _22545_/X _22548_/X _22549_/X _22550_/X vssd1 vssd1 vccd1
+ vccd1 _22556_/A sky130_fd_sc_hd__mux4_1
XFILLER_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21506_ _21506_/A vssd1 vssd1 vccd1 vccd1 _21506_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25274_ _25306_/A _25274_/B vssd1 vssd1 vccd1 vccd1 _25274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_195_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22486_ _22486_/A vssd1 vssd1 vccd1 vccd1 _22486_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27013_ _22850_/X _27013_/D vssd1 vssd1 vccd1 vccd1 _27013_/Q sky130_fd_sc_hd__dfxtp_1
X_24225_ _24225_/A _24235_/B vssd1 vssd1 vccd1 vccd1 _27382_/D sky130_fd_sc_hd__nor2_1
X_21437_ _21427_/X _21428_/X _21429_/X _21430_/X _21431_/X _21432_/X vssd1 vssd1 vccd1
+ vccd1 _21438_/A sky130_fd_sc_hd__mux4_1
XFILLER_182_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24156_ _27455_/Q _24162_/B vssd1 vssd1 vccd1 vccd1 _24157_/A sky130_fd_sc_hd__and2_1
X_21368_ _21368_/A vssd1 vssd1 vccd1 vccd1 _21368_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23107_ _27097_/Q _17775_/X _23107_/S vssd1 vssd1 vccd1 vccd1 _23108_/A sky130_fd_sc_hd__mux2_1
X_20319_ _20335_/A vssd1 vssd1 vccd1 vccd1 _20319_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24087_ _27392_/Q _24095_/B vssd1 vssd1 vccd1 vccd1 _24088_/A sky130_fd_sc_hd__and2_1
X_21299_ _21285_/X _21286_/X _21287_/X _21288_/X _21289_/X _21290_/X vssd1 vssd1 vccd1
+ vccd1 _21300_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23038_ _23094_/A vssd1 vssd1 vccd1 vccd1 _23107_/S sky130_fd_sc_hd__buf_2
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_472 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27846_ _27850_/CLK _27846_/D vssd1 vssd1 vccd1 vccd1 _27846_/Q sky130_fd_sc_hd__dfxtp_1
X_15860_ _15862_/A vssd1 vssd1 vccd1 vccd1 _15860_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14811_ _14810_/X _26522_/Q _14811_/S vssd1 vssd1 vccd1 vccd1 _14812_/A sky130_fd_sc_hd__mux2_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27777_ _27784_/CLK _27777_/D vssd1 vssd1 vccd1 vccd1 _27777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15791_ _15791_/A vssd1 vssd1 vccd1 vccd1 _26103_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24989_ _27964_/A _24987_/X _25024_/S vssd1 vssd1 vccd1 vccd1 _24990_/A sky130_fd_sc_hd__mux2_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _17586_/A vssd1 vssd1 vccd1 vccd1 _17599_/S sky130_fd_sc_hd__buf_2
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26728_ _21860_/X _26728_/D vssd1 vssd1 vccd1 vccd1 _26728_/Q sky130_fd_sc_hd__dfxtp_1
X_14742_ _14742_/A vssd1 vssd1 vccd1 vccd1 _26544_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14673_ _26568_/Q _14671_/X _14666_/X _14672_/Y vssd1 vssd1 vccd1 vccd1 _26568_/D
+ sky130_fd_sc_hd__a31o_1
X_17461_ _17460_/X _25822_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17462_/A sky130_fd_sc_hd__mux2_1
X_26659_ _21614_/X _26659_/D vssd1 vssd1 vccd1 vccd1 _26659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19200_ _19190_/X _19195_/X _19199_/X _19151_/X _19105_/X vssd1 vssd1 vccd1 vccd1
+ _19201_/C sky130_fd_sc_hd__a221o_1
X_13624_ _13895_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16412_ _16412_/A vssd1 vssd1 vccd1 vccd1 _16412_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17392_ input6/X vssd1 vssd1 vccd1 vccd1 _20792_/A sky130_fd_sc_hd__inv_2
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19131_ _19131_/A vssd1 vssd1 vccd1 vccd1 _26053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13555_ _14511_/A vssd1 vssd1 vccd1 vccd1 _13926_/A sky130_fd_sc_hd__buf_2
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16343_ _14807_/A _16384_/A _16374_/A _25945_/Q _16342_/Y vssd1 vssd1 vccd1 vccd1
+ _16862_/B sky130_fd_sc_hd__a221o_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater77 _27430_/CLK vssd1 vssd1 vccd1 vccd1 _27436_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater88 _27219_/CLK vssd1 vssd1 vccd1 vccd1 _27422_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_13_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater99 _27219_/CLK vssd1 vssd1 vccd1 vccd1 _27294_/CLK sky130_fd_sc_hd__clkbuf_1
X_19062_ _26947_/Q _26915_/Q _26883_/Q _26851_/Q _19061_/X _18898_/X vssd1 vssd1 vccd1
+ vccd1 _19062_/X sky130_fd_sc_hd__mux4_2
X_16274_ _26060_/Q _16274_/B _16274_/C vssd1 vssd1 vccd1 vccd1 _16274_/X sky130_fd_sc_hd__and3_1
X_13486_ _26959_/Q _13464_/X _13482_/X _13485_/Y vssd1 vssd1 vccd1 vccd1 _26959_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18013_ _26816_/Q _26784_/Q _26752_/Q _26720_/Q _18011_/X _24388_/A vssd1 vssd1 vccd1
+ vccd1 _18013_/X sky130_fd_sc_hd__mux4_1
X_15225_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15234_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15156_ _26377_/Q _13373_/X _15162_/S vssd1 vssd1 vccd1 vccd1 _15157_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14107_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15087_ _15087_/A vssd1 vssd1 vccd1 vccd1 _26408_/D sky130_fd_sc_hd__clkbuf_1
X_19964_ _19956_/X _19957_/X _19958_/X _19959_/X _19960_/X _19961_/X vssd1 vssd1 vccd1
+ vccd1 _19965_/A sky130_fd_sc_hd__mux4_1
X_18915_ _18930_/A vssd1 vssd1 vccd1 vccd1 _24400_/A sky130_fd_sc_hd__buf_4
X_14038_ _14038_/A vssd1 vssd1 vccd1 vccd1 _14038_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19895_ _19895_/A vssd1 vssd1 vccd1 vccd1 _19895_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18846_ _18969_/A _18846_/B vssd1 vssd1 vccd1 vccd1 _18846_/X sky130_fd_sc_hd__or2_1
XFILLER_41_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_518 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18777_ _18922_/A vssd1 vssd1 vccd1 vccd1 _18913_/A sky130_fd_sc_hd__clkbuf_4
X_15989_ _27753_/Q vssd1 vssd1 vccd1 vccd1 _25430_/A sky130_fd_sc_hd__inv_2
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17728_ _27424_/Q vssd1 vssd1 vccd1 vccd1 _17728_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17659_ _17504_/X _25900_/Q _17667_/S vssd1 vssd1 vccd1 vccd1 _17660_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20670_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19329_ _26286_/Q _26254_/Q _26222_/Q _26190_/Q _19283_/X _19192_/X vssd1 vssd1 vccd1
+ vccd1 _19329_/X sky130_fd_sc_hd__mux4_1
XFILLER_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22340_ _22340_/A vssd1 vssd1 vccd1 vccd1 _22340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22271_ _22261_/X _22262_/X _22263_/X _22264_/X _22266_/X _22268_/X vssd1 vssd1 vccd1
+ vccd1 _22272_/A sky130_fd_sc_hd__mux4_1
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24010_ _27092_/Q _27124_/Q _24032_/S vssd1 vssd1 vccd1 vccd1 _24010_/X sky130_fd_sc_hd__mux2_1
X_21222_ _21222_/A vssd1 vssd1 vccd1 vccd1 _21222_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21153_ _21144_/X _21146_/X _21148_/X _21150_/X _21151_/X _21152_/X vssd1 vssd1 vccd1
+ vccd1 _21154_/A sky130_fd_sc_hd__mux4_1
XFILLER_137_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20104_ _20095_/X _20097_/X _20099_/X _20101_/X _20102_/X _20103_/X vssd1 vssd1 vccd1
+ vccd1 _20105_/A sky130_fd_sc_hd__mux4_1
XFILLER_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21084_ _21084_/A vssd1 vssd1 vccd1 vccd1 _21084_/X sky130_fd_sc_hd__clkbuf_1
X_25961_ _25963_/CLK _25961_/D vssd1 vssd1 vccd1 vccd1 _25961_/Q sky130_fd_sc_hd__dfxtp_1
X_27700_ _27700_/CLK _27700_/D vssd1 vssd1 vccd1 vccd1 _27700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24912_ _24918_/B _24912_/B vssd1 vssd1 vccd1 vccd1 _24913_/B sky130_fd_sc_hd__or2_1
X_20035_ _20035_/A vssd1 vssd1 vccd1 vccd1 _20035_/X sky130_fd_sc_hd__clkbuf_1
X_25892_ _25941_/CLK _25892_/D vssd1 vssd1 vccd1 vccd1 _25892_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27631_ _27633_/CLK _27631_/D vssd1 vssd1 vccd1 vccd1 _27631_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24843_ _27758_/Q _27757_/Q _27756_/Q _27755_/Q vssd1 vssd1 vccd1 vccd1 _24851_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24774_ _27623_/Q _24771_/X _24772_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _27623_/D
+ sky130_fd_sc_hd__o211a_1
X_27562_ _27562_/CLK _27562_/D vssd1 vssd1 vccd1 vccd1 _27562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _21986_/A vssd1 vssd1 vccd1 vccd1 _21986_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26513_ _21106_/X _26513_/D vssd1 vssd1 vccd1 vccd1 _26513_/Q sky130_fd_sc_hd__dfxtp_1
X_23725_ _27369_/Q _24005_/A vssd1 vssd1 vccd1 vccd1 _23726_/A sky130_fd_sc_hd__and2_1
X_20937_ _20953_/A vssd1 vssd1 vccd1 vccd1 _20937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27493_ _27495_/CLK _27493_/D vssd1 vssd1 vccd1 vccd1 _27493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26444_ _20863_/X _26444_/D vssd1 vssd1 vccd1 vccd1 _26444_/Q sky130_fd_sc_hd__dfxtp_1
X_23656_ _23656_/A vssd1 vssd1 vccd1 vccd1 _27234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _25639_/A vssd1 vssd1 vccd1 vccd1 _21215_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22607_ _22593_/X _22594_/X _22595_/X _22596_/X _22597_/X _22598_/X vssd1 vssd1 vccd1
+ vccd1 _22608_/A sky130_fd_sc_hd__mux4_1
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26375_ _20627_/X _26375_/D vssd1 vssd1 vccd1 vccd1 _26375_/Q sky130_fd_sc_hd__dfxtp_1
X_23587_ _23587_/A vssd1 vssd1 vccd1 vccd1 _27216_/D sky130_fd_sc_hd__clkbuf_1
X_20799_ _20866_/A vssd1 vssd1 vccd1 vccd1 _20799_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25326_ _25344_/A _25326_/B vssd1 vssd1 vccd1 vccd1 _25326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ _13340_/A vssd1 vssd1 vccd1 vccd1 _26996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22538_ _22887_/A vssd1 vssd1 vccd1 vccd1 _22609_/A sky130_fd_sc_hd__buf_2
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25257_ _27538_/Q _27506_/Q vssd1 vssd1 vccd1 vccd1 _25258_/B sky130_fd_sc_hd__and2_1
XFILLER_5_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13271_ _13317_/S vssd1 vssd1 vccd1 vccd1 _13280_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22469_ _22452_/X _22454_/X _22456_/X _22458_/X _22459_/X _22460_/X vssd1 vssd1 vccd1
+ vccd1 _22470_/A sky130_fd_sc_hd__mux4_1
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15010_ _15023_/A vssd1 vssd1 vccd1 vccd1 _15021_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24208_ _24208_/A _24210_/B vssd1 vssd1 vccd1 vccd1 _27372_/D sky130_fd_sc_hd__nor2_1
XFILLER_170_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25188_ _25188_/A _25187_/X vssd1 vssd1 vccd1 vccd1 _25191_/A sky130_fd_sc_hd__or2b_1
XFILLER_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24139_ _24139_/A vssd1 vssd1 vccd1 vccd1 _27342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_842 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16961_ _27590_/Q vssd1 vssd1 vccd1 vccd1 _16971_/B sky130_fd_sc_hd__inv_2
X_18700_ _26013_/Q _17686_/X _18702_/S vssd1 vssd1 vccd1 vccd1 _18701_/A sky130_fd_sc_hd__mux2_1
X_15912_ _15912_/A vssd1 vssd1 vccd1 vccd1 _15912_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19680_ _19728_/A vssd1 vssd1 vccd1 vccd1 _19680_/X sky130_fd_sc_hd__clkbuf_1
X_16892_ _16077_/A _16772_/A _16479_/A _16621_/X vssd1 vssd1 vccd1 vccd1 _16892_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18631_ _18631_/A vssd1 vssd1 vccd1 vccd1 _25982_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _13210_/X _26079_/Q _15849_/S vssd1 vssd1 vccd1 vccd1 _15844_/A sky130_fd_sc_hd__mux2_1
X_27829_ _27830_/CLK _27829_/D vssd1 vssd1 vccd1 vccd1 _27829_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18562_ _18560_/X _18561_/X _18580_/S vssd1 vssd1 vccd1 vccd1 _18562_/X sky130_fd_sc_hd__mux2_2
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _23562_/A vssd1 vssd1 vccd1 vccd1 _15774_/X sky130_fd_sc_hd__clkbuf_4
X_12986_ _12986_/A vssd1 vssd1 vccd1 vccd1 _27805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17513_ _17513_/A vssd1 vssd1 vccd1 vccd1 _25838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14725_ _14724_/X _26549_/Q _14725_/S vssd1 vssd1 vccd1 vccd1 _14726_/A sky130_fd_sc_hd__mux2_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _27820_/Q _26581_/Q _26453_/Q _26133_/Q _18401_/X _18425_/X vssd1 vssd1 vccd1
+ vccd1 _18493_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _27414_/Q vssd1 vssd1 vccd1 vccd1 _17444_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14656_ _15730_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14656_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13607_ _26931_/Q _13599_/X _13603_/X _13606_/Y vssd1 vssd1 vccd1 vccd1 _26931_/D
+ sky130_fd_sc_hd__a31o_1
X_17375_ _27096_/Q _27128_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17375_/X sky130_fd_sc_hd__mux2_1
X_14587_ _15749_/A _14597_/B vssd1 vssd1 vccd1 vccd1 _14587_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19114_ _26693_/Q _26661_/Q _26629_/Q _26597_/Q _19015_/X _19087_/X vssd1 vssd1 vccd1
+ vccd1 _19114_/X sky130_fd_sc_hd__mux4_2
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16326_ _16326_/A vssd1 vssd1 vccd1 vccd1 _16752_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_1030 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13538_ _13915_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19045_ _26946_/Q _26914_/Q _26882_/Q _26850_/Q _19044_/X _18972_/X vssd1 vssd1 vccd1
+ vccd1 _19045_/X sky130_fd_sc_hd__mux4_2
X_16257_ _16257_/A vssd1 vssd1 vccd1 vccd1 _16292_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13469_ _27359_/Q _13108_/X _13029_/A _27327_/Q _13097_/X vssd1 vssd1 vccd1 vccd1
+ _16563_/A sky130_fd_sc_hd__a221oi_4
XFILLER_173_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15208_ _14734_/X _26354_/Q _15212_/S vssd1 vssd1 vccd1 vccd1 _15209_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16188_ _26044_/Q _16191_/B _16194_/C vssd1 vssd1 vccd1 vccd1 _16188_/X sky130_fd_sc_hd__and3_1
XFILLER_182_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _15139_/A vssd1 vssd1 vccd1 vccd1 _26385_/D sky130_fd_sc_hd__clkbuf_1
X_19947_ _19947_/A vssd1 vssd1 vccd1 vccd1 _19947_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ _19866_/X _19867_/X _19868_/X _19869_/X _19870_/X _19871_/X vssd1 vssd1 vccd1
+ vccd1 _19879_/A sky130_fd_sc_hd__mux4_1
XFILLER_96_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18829_ _19414_/A vssd1 vssd1 vccd1 vccd1 _18829_/X sky130_fd_sc_hd__buf_4
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21840_ _21840_/A vssd1 vssd1 vccd1 vccd1 _21840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21771_ _21758_/X _21760_/X _21762_/X _21764_/X _21765_/X _21766_/X vssd1 vssd1 vccd1
+ vccd1 _21772_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23510_ _25976_/Q _27195_/Q _23525_/S vssd1 vssd1 vccd1 vccd1 _23511_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20722_ _20770_/A vssd1 vssd1 vccd1 vccd1 _20722_/X sky130_fd_sc_hd__clkbuf_1
X_24490_ _27584_/Q _27583_/Q _27579_/Q _27578_/Q vssd1 vssd1 vccd1 vccd1 _24491_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_196_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23441_ input39/X _23429_/X _23440_/X _23434_/X vssd1 vssd1 vccd1 vccd1 _27170_/D
+ sky130_fd_sc_hd__o211a_1
X_20653_ _20685_/A vssd1 vssd1 vccd1 vccd1 _20653_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26160_ _19873_/X _26160_/D vssd1 vssd1 vccd1 vccd1 _26160_/Q sky130_fd_sc_hd__dfxtp_1
X_23372_ _24778_/A _27250_/Q _27251_/Q _24780_/A vssd1 vssd1 vccd1 vccd1 _23372_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_20584_ _20600_/A vssd1 vssd1 vccd1 vccd1 _20584_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25111_ _25143_/A vssd1 vssd1 vccd1 vccd1 _25356_/A sky130_fd_sc_hd__clkbuf_2
X_22323_ _22315_/X _22316_/X _22317_/X _22318_/X _22319_/X _22320_/X vssd1 vssd1 vccd1
+ vccd1 _22324_/A sky130_fd_sc_hd__mux4_1
X_26091_ _19630_/X _26091_/D vssd1 vssd1 vccd1 vccd1 _26091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25042_ _27970_/A _25041_/X _25067_/S vssd1 vssd1 vccd1 vccd1 _25043_/A sky130_fd_sc_hd__mux2_1
X_22254_ _22254_/A vssd1 vssd1 vccd1 vccd1 _22254_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21205_ _21195_/X _21196_/X _21197_/X _21198_/X _21199_/X _21200_/X vssd1 vssd1 vccd1
+ vccd1 _21206_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22185_ _22173_/X _22174_/X _22175_/X _22176_/X _22179_/X _22182_/X vssd1 vssd1 vccd1
+ vccd1 _22186_/A sky130_fd_sc_hd__mux4_1
XFILLER_133_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21136_ _21136_/A vssd1 vssd1 vccd1 vccd1 _21136_/X sky130_fd_sc_hd__clkbuf_1
X_26993_ _22780_/X _26993_/D vssd1 vssd1 vccd1 vccd1 _26993_/Q sky130_fd_sc_hd__dfxtp_1
X_21067_ _21058_/X _21060_/X _21062_/X _21064_/X _21065_/X _21066_/X vssd1 vssd1 vccd1
+ vccd1 _21068_/A sky130_fd_sc_hd__mux4_1
X_25944_ _26047_/CLK _25944_/D vssd1 vssd1 vccd1 vccd1 _25944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20018_ _20009_/X _20011_/X _20013_/X _20015_/X _20016_/X _20017_/X vssd1 vssd1 vccd1
+ vccd1 _20019_/A sky130_fd_sc_hd__mux4_2
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25875_ _27130_/CLK _25875_/D vssd1 vssd1 vccd1 vccd1 _25875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27614_ _27614_/CLK _27614_/D vssd1 vssd1 vccd1 vccd1 _27614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24826_ _27641_/Q _24813_/X _24825_/Y _24817_/X vssd1 vssd1 vccd1 vccd1 _27641_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27545_ _27564_/CLK _27545_/D vssd1 vssd1 vccd1 vccd1 _27545_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21969_ _21985_/A vssd1 vssd1 vccd1 vccd1 _21969_/X sky130_fd_sc_hd__clkbuf_2
X_24757_ _27617_/Q _24742_/X _24756_/Y _24746_/X vssd1 vssd1 vccd1 vccd1 _27617_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _14510_/A vssd1 vssd1 vccd1 vccd1 _14510_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23708_ _24941_/A _27258_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23709_/A sky130_fd_sc_hd__mux2_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _13078_/X _26229_/Q _15490_/S vssd1 vssd1 vccd1 vccd1 _15491_/A sky130_fd_sc_hd__mux2_1
X_24688_ _25540_/A vssd1 vssd1 vccd1 vccd1 _24698_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27476_ _27477_/CLK _27476_/D vssd1 vssd1 vccd1 vccd1 _27476_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14441_ _14441_/A vssd1 vssd1 vccd1 vccd1 _14441_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26427_ _20811_/X _26427_/D vssd1 vssd1 vccd1 vccd1 _26427_/Q sky130_fd_sc_hd__dfxtp_1
X_23639_ _23638_/A _27227_/Q _27228_/Q _23638_/B vssd1 vssd1 vccd1 vccd1 _23640_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14372_ _14372_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14372_/Y sky130_fd_sc_hd__nor2_1
X_17160_ _17120_/X _17158_/X _17159_/X vssd1 vssd1 vccd1 vccd1 _17160_/X sky130_fd_sc_hd__a21bo_1
XFILLER_122_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26358_ _20563_/X _26358_/D vssd1 vssd1 vccd1 vccd1 _26358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _26072_/Q vssd1 vssd1 vccd1 vccd1 _16111_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ _27001_/Q _13319_/X _13335_/S vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__mux2_1
X_25309_ _25309_/A vssd1 vssd1 vccd1 vccd1 _25344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26289_ _20317_/X _26289_/D vssd1 vssd1 vccd1 vccd1 _26289_/Q sky130_fd_sc_hd__dfxtp_1
X_17091_ _27201_/Q _17090_/X _17128_/S vssd1 vssd1 vccd1 vccd1 _17092_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16042_ _16062_/A _16062_/B _16040_/Y _16041_/X vssd1 vssd1 vccd1 vccd1 _16066_/A
+ sky130_fd_sc_hd__o211a_1
X_13254_ _27031_/Q _13067_/X _13258_/S vssd1 vssd1 vccd1 vccd1 _13255_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ _27043_/Q _13184_/X _13199_/S vssd1 vssd1 vccd1 vccd1 _13186_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19801_ _19801_/A vssd1 vssd1 vccd1 vccd1 _19801_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ _17993_/A vssd1 vssd1 vccd1 vccd1 _25949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19732_ _25726_/A vssd1 vssd1 vccd1 vccd1 _19801_/A sky130_fd_sc_hd__clkbuf_2
X_16944_ _27600_/Q _24208_/A _24206_/A _27598_/Q _16943_/X vssd1 vssd1 vccd1 vccd1
+ _16945_/C sky130_fd_sc_hd__o221a_1
XFILLER_1_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19663_ _19728_/A vssd1 vssd1 vccd1 vccd1 _19663_/X sky130_fd_sc_hd__clkbuf_1
X_16875_ _24226_/A _24235_/A _24237_/A _16875_/D vssd1 vssd1 vccd1 vccd1 _16875_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18614_ _25568_/A _25115_/A vssd1 vssd1 vccd1 vccd1 _18614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _15826_/A vssd1 vssd1 vccd1 vccd1 _26087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19594_ _19626_/A vssd1 vssd1 vccd1 vccd1 _19594_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18545_ _18539_/X _18541_/X _18544_/X _18443_/X _18489_/X vssd1 vssd1 vccd1 vccd1
+ _18546_/C sky130_fd_sc_hd__a221o_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _26116_/Q _15747_/X _15753_/X _15756_/Y vssd1 vssd1 vccd1 vccd1 _26116_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _12969_/A vssd1 vssd1 vccd1 vccd1 _27813_/D sky130_fd_sc_hd__clkbuf_1
X_14708_ _26554_/Q _14698_/X _14631_/B _14707_/Y vssd1 vssd1 vccd1 vccd1 _26554_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_61_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18476_ _18379_/X _18472_/X _18475_/X _18384_/X vssd1 vssd1 vccd1 vccd1 _18476_/X
+ sky130_fd_sc_hd__o211a_1
X_15688_ _15688_/A vssd1 vssd1 vccd1 vccd1 _26141_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_380 _15773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17427_ _17427_/A vssd1 vssd1 vccd1 vccd1 _25811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14639_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17358_ _17358_/A vssd1 vssd1 vccd1 vccd1 _27944_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_159_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16309_ _16309_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16309_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ _25935_/Q _26001_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17290_/B sky130_fd_sc_hd__mux2_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19028_ _19441_/A vssd1 vssd1 vccd1 vccd1 _19028_/X sky130_fd_sc_hd__buf_2
XFILLER_177_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23990_ _23990_/A vssd1 vssd1 vccd1 vccd1 _23990_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_559 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22941_ _22957_/A vssd1 vssd1 vccd1 vccd1 _22941_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22872_ _22872_/A vssd1 vssd1 vccd1 vccd1 _22872_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25660_ _25724_/A vssd1 vssd1 vccd1 vccd1 _25660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21823_ _21809_/X _21810_/X _21811_/X _21812_/X _21813_/X _21814_/X vssd1 vssd1 vccd1
+ vccd1 _21824_/A sky130_fd_sc_hd__mux4_1
X_24611_ _24611_/A vssd1 vssd1 vccd1 vccd1 _24620_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_83_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25591_ _27715_/Q _25433_/X _25435_/X vssd1 vssd1 vccd1 vccd1 _25591_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27330_ _27402_/CLK _27330_/D vssd1 vssd1 vccd1 vccd1 _27330_/Q sky130_fd_sc_hd__dfxtp_1
X_24542_ _24534_/X _24388_/A _24545_/S vssd1 vssd1 vccd1 vccd1 _24543_/B sky130_fd_sc_hd__mux2_1
X_21754_ _21754_/A vssd1 vssd1 vccd1 vccd1 _21754_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20705_ _20771_/A vssd1 vssd1 vccd1 vccd1 _20705_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24473_ _24473_/A vssd1 vssd1 vccd1 vccd1 _27512_/D sky130_fd_sc_hd__clkbuf_1
X_27261_ _27261_/CLK _27261_/D vssd1 vssd1 vccd1 vccd1 _27261_/Q sky130_fd_sc_hd__dfxtp_1
X_21685_ _21667_/X _21670_/X _21673_/X _21676_/X _21677_/X _21678_/X vssd1 vssd1 vccd1
+ vccd1 _21686_/A sky130_fd_sc_hd__mux4_1
XFILLER_196_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26212_ _20055_/X _26212_/D vssd1 vssd1 vccd1 vccd1 _26212_/Q sky130_fd_sc_hd__dfxtp_1
X_23424_ input20/X _23415_/X _23423_/X _23421_/X vssd1 vssd1 vccd1 vccd1 _27163_/D
+ sky130_fd_sc_hd__o211a_1
X_27192_ _27536_/CLK _27192_/D vssd1 vssd1 vccd1 vccd1 _27192_/Q sky130_fd_sc_hd__dfxtp_1
X_20636_ _20684_/A vssd1 vssd1 vccd1 vccd1 _20636_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26143_ _19809_/X _26143_/D vssd1 vssd1 vccd1 vccd1 _26143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23355_ _27781_/Q vssd1 vssd1 vccd1 vccd1 _24808_/A sky130_fd_sc_hd__inv_2
X_20567_ _20599_/A vssd1 vssd1 vccd1 vccd1 _20567_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22306_ _22306_/A vssd1 vssd1 vccd1 vccd1 _22306_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26074_ _17407_/A _26074_/D vssd1 vssd1 vccd1 vccd1 _26074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23286_ _27752_/Q input65/X vssd1 vssd1 vccd1 vccd1 _23286_/X sky130_fd_sc_hd__xor2_1
X_20498_ _20514_/A vssd1 vssd1 vccd1 vccd1 _20498_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25025_ _25025_/A vssd1 vssd1 vccd1 vccd1 _27677_/D sky130_fd_sc_hd__clkbuf_1
X_22237_ _22229_/X _22230_/X _22231_/X _22232_/X _22233_/X _22234_/X vssd1 vssd1 vccd1
+ vccd1 _22238_/A sky130_fd_sc_hd__mux4_1
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22168_ _22168_/A vssd1 vssd1 vccd1 vccd1 _22168_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21119_ _21109_/X _21110_/X _21111_/X _21112_/X _21113_/X _21114_/X vssd1 vssd1 vccd1
+ vccd1 _21120_/A sky130_fd_sc_hd__mux4_1
XFILLER_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22099_ _22083_/X _22084_/X _22085_/X _22086_/X _22088_/X _22090_/X vssd1 vssd1 vccd1
+ vccd1 _22100_/A sky130_fd_sc_hd__mux4_1
X_14990_ _15728_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14990_/Y sky130_fd_sc_hd__nor2_1
X_26976_ _22728_/X _26976_/D vssd1 vssd1 vccd1 vccd1 _26976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _26810_/Q _13933_/X _13861_/B _13940_/Y vssd1 vssd1 vccd1 vccd1 _26810_/D
+ sky130_fd_sc_hd__a31o_1
X_25927_ _27144_/CLK _25927_/D vssd1 vssd1 vccd1 vccd1 _25927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16660_ _16660_/A _16885_/A vssd1 vssd1 vccd1 vccd1 _16660_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13872_ _13872_/A vssd1 vssd1 vccd1 vccd1 _13925_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_25858_ _27842_/CLK _25858_/D vssd1 vssd1 vccd1 vccd1 _25858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15611_ _26175_/Q _16224_/A _15617_/S vssd1 vssd1 vccd1 vccd1 _15612_/A sky130_fd_sc_hd__mux2_1
X_24809_ _27636_/Q _24798_/X _24808_/Y _24801_/X vssd1 vssd1 vccd1 vccd1 _27636_/D
+ sky130_fd_sc_hd__o211a_1
X_16591_ _25972_/Q _16098_/X _16590_/X vssd1 vssd1 vccd1 vccd1 _16791_/B sky130_fd_sc_hd__a21oi_2
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25789_ _25789_/A vssd1 vssd1 vccd1 vccd1 _27849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18330_ _26413_/Q _26381_/Q _26349_/Q _26317_/Q _18305_/X _18329_/X vssd1 vssd1 vccd1
+ vccd1 _18330_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27528_ _27604_/CLK _27528_/D vssd1 vssd1 vccd1 vccd1 _27528_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _15542_/A vssd1 vssd1 vccd1 vccd1 _26206_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18261_ _26410_/Q _26378_/Q _26346_/Q _26314_/Q _18189_/X _18214_/X vssd1 vssd1 vccd1
+ vccd1 _18261_/X sky130_fd_sc_hd__mux4_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27459_ _27462_/CLK _27459_/D vssd1 vssd1 vccd1 vccd1 _27459_/Q sky130_fd_sc_hd__dfxtp_1
X_15473_ _26236_/Q _13414_/X _15473_/S vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17210_/X _17211_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17212_/X sky130_fd_sc_hd__mux2_1
X_14424_ _26648_/Q _14421_/X _14416_/X _14423_/Y vssd1 vssd1 vccd1 vccd1 _26648_/D
+ sky130_fd_sc_hd__a31o_1
X_18192_ _18184_/X _18187_/X _18191_/X _18168_/X _18122_/X vssd1 vssd1 vccd1 vccd1
+ _18193_/C sky130_fd_sc_hd__a221o_1
XFILLER_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ _27837_/Q _27141_/Q _25886_/Q _25854_/Q _17142_/X _17130_/X vssd1 vssd1 vccd1
+ vccd1 _17143_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14355_ _26673_/Q _14352_/X _14345_/X _14354_/Y vssd1 vssd1 vccd1 vccd1 _26673_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13306_ _13306_/A vssd1 vssd1 vccd1 vccd1 _27008_/D sky130_fd_sc_hd__clkbuf_1
X_14286_ _26698_/Q _14283_/X _14284_/X _14285_/Y vssd1 vssd1 vccd1 vccd1 _26698_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17074_ _17057_/X _17073_/X _17033_/X vssd1 vssd1 vccd1 vccd1 _17074_/X sky130_fd_sc_hd__a21bo_1
XFILLER_170_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ _27271_/Q _13237_/B vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__and2_1
X_16025_ _16252_/C vssd1 vssd1 vccd1 vccd1 _16296_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ _13168_/A vssd1 vssd1 vccd1 vccd1 _27046_/D sky130_fd_sc_hd__clkbuf_1
X_17976_ _26815_/Q _26783_/Q _26751_/Q _26719_/Q _17863_/X _17890_/X vssd1 vssd1 vccd1
+ vccd1 _17976_/X sky130_fd_sc_hd__mux4_1
X_13099_ _14734_/A vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__buf_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19715_ _19715_/A vssd1 vssd1 vccd1 vccd1 _19715_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16927_ _27594_/Q _24207_/A _24206_/A _27593_/Q vssd1 vssd1 vccd1 vccd1 _16927_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19646_ _25726_/A vssd1 vssd1 vccd1 vccd1 _19715_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16858_ _16858_/A _16858_/B vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_81_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15809_ _15809_/A vssd1 vssd1 vccd1 vccd1 _26095_/D sky130_fd_sc_hd__clkbuf_1
X_19577_ _19625_/A vssd1 vssd1 vccd1 vccd1 _19577_/X sky130_fd_sc_hd__clkbuf_2
X_16789_ _16110_/A _24309_/A _16559_/A vssd1 vssd1 vccd1 vccd1 _16790_/B sky130_fd_sc_hd__o21ai_2
XFILLER_81_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18528_ _18842_/A _18528_/B _18528_/C vssd1 vssd1 vccd1 vccd1 _18529_/A sky130_fd_sc_hd__and3_1
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18459_ _26291_/Q _26259_/Q _26227_/Q _26195_/Q _18458_/X _18324_/X vssd1 vssd1 vccd1
+ vccd1 _18459_/X sky130_fd_sc_hd__mux4_1
X_27960__446 vssd1 vssd1 vccd1 vccd1 _27960__446/HI _27960_/A sky130_fd_sc_hd__conb_1
X_21470_ _21470_/A vssd1 vssd1 vccd1 vccd1 _21470_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20421_ _20421_/A vssd1 vssd1 vccd1 vccd1 _20421_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23140_ _23140_/A vssd1 vssd1 vccd1 vccd1 _27110_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20352_ _25653_/A vssd1 vssd1 vccd1 vccd1 _20702_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23071_ _23071_/A vssd1 vssd1 vccd1 vccd1 _27080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20283_ _20283_/A vssd1 vssd1 vccd1 vccd1 _20283_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22022_ _22086_/A vssd1 vssd1 vccd1 vccd1 _22022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26830_ _22220_/X _26830_/D vssd1 vssd1 vccd1 vccd1 _26830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26761_ _21974_/X _26761_/D vssd1 vssd1 vccd1 vccd1 _26761_/Q sky130_fd_sc_hd__dfxtp_1
X_23973_ _27088_/Q _23954_/X _23955_/X _27120_/Q _23956_/X vssd1 vssd1 vccd1 vccd1
+ _23973_/X sky130_fd_sc_hd__a221o_1
XFILLER_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25712_ _25712_/A vssd1 vssd1 vccd1 vccd1 _25712_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22924_ _22956_/A vssd1 vssd1 vccd1 vccd1 _22924_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26692_ _21732_/X _26692_/D vssd1 vssd1 vccd1 vccd1 _26692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25643_ _25635_/X _25636_/X _25637_/X _25638_/X _25640_/X _25642_/X vssd1 vssd1 vccd1
+ vccd1 _25644_/A sky130_fd_sc_hd__mux4_1
X_22855_ _22871_/A vssd1 vssd1 vccd1 vccd1 _22855_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21806_ _21806_/A vssd1 vssd1 vccd1 vccd1 _21806_/X sky130_fd_sc_hd__clkbuf_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25574_ _25560_/X _25296_/B _25573_/X _25566_/X vssd1 vssd1 vccd1 vccd1 _25574_/X
+ sky130_fd_sc_hd__a211o_1
X_22786_ _22786_/A vssd1 vssd1 vccd1 vccd1 _22786_/X sky130_fd_sc_hd__clkbuf_1
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27313_ _27334_/CLK _27313_/D vssd1 vssd1 vccd1 vccd1 _27313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21737_ _21737_/A vssd1 vssd1 vccd1 vccd1 _21737_/X sky130_fd_sc_hd__clkbuf_1
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24525_ _27585_/Q _24633_/A _24522_/A _24631_/B _24398_/A vssd1 vssd1 vccd1 vccd1
+ _24525_/X sky130_fd_sc_hd__a32o_1
XFILLER_200_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27244_ _27262_/CLK _27244_/D vssd1 vssd1 vccd1 vccd1 _27244_/Q sky130_fd_sc_hd__dfxtp_1
X_21668_ _22540_/A vssd1 vssd1 vccd1 vccd1 _22017_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24456_ _27626_/Q _24456_/B vssd1 vssd1 vccd1 vccd1 _24457_/A sky130_fd_sc_hd__and2_1
XFILLER_71_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20619_ _20685_/A vssd1 vssd1 vccd1 vccd1 _20619_/X sky130_fd_sc_hd__clkbuf_1
X_23407_ _24823_/A _27233_/Q _27239_/Q _24750_/A vssd1 vssd1 vccd1 vccd1 _23407_/X
+ sky130_fd_sc_hd__o22a_1
X_27175_ _27608_/CLK _27175_/D vssd1 vssd1 vccd1 vccd1 _27175_/Q sky130_fd_sc_hd__dfxtp_1
X_24387_ _24387_/A vssd1 vssd1 vccd1 vccd1 _27474_/D sky130_fd_sc_hd__clkbuf_1
X_21599_ _21647_/A vssd1 vssd1 vccd1 vccd1 _21599_/X sky130_fd_sc_hd__clkbuf_1
X_14140_ _14406_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _14140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26126_ _19757_/X _26126_/D vssd1 vssd1 vccd1 vccd1 _26126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23338_ _27777_/Q vssd1 vssd1 vccd1 vccd1 _24796_/A sky130_fd_sc_hd__inv_2
XFILLER_138_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14071_ _26775_/Q _14058_/X _14064_/X _14070_/Y vssd1 vssd1 vccd1 vccd1 _26775_/D
+ sky130_fd_sc_hd__a31o_1
X_23269_ _27734_/Q _23267_/Y _23268_/Y input58/X vssd1 vssd1 vccd1 vccd1 _23269_/X
+ sky130_fd_sc_hd__o22a_1
X_26057_ _26057_/CLK _26057_/D vssd1 vssd1 vccd1 vccd1 _26057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13022_ _13529_/A vssd1 vssd1 vccd1 vccd1 _13022_/X sky130_fd_sc_hd__clkbuf_4
X_25008_ _27830_/Q _27134_/Q _25879_/Q _25847_/Q _24972_/X _24991_/X vssd1 vssd1 vccd1
+ vccd1 _25008_/X sky130_fd_sc_hd__mux4_1
XFILLER_105_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17830_ _18020_/A vssd1 vssd1 vccd1 vccd1 _17830_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17761_ _25938_/Q _17760_/X _17770_/S vssd1 vssd1 vccd1 vccd1 _17762_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26959_ _22664_/X _26959_/D vssd1 vssd1 vccd1 vccd1 _26959_/Q sky130_fd_sc_hd__dfxtp_1
X_14973_ _26453_/Q _14957_/X _14960_/X _14972_/Y vssd1 vssd1 vccd1 vccd1 _26453_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19500_ _26710_/Q _26678_/Q _26646_/Q _26614_/Q _18767_/X _18909_/X vssd1 vssd1 vccd1
+ vccd1 _19501_/B sky130_fd_sc_hd__mux4_1
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16712_ _16625_/A _16774_/A _16711_/Y _16625_/B vssd1 vssd1 vccd1 vccd1 _16712_/X
+ sky130_fd_sc_hd__a31o_1
X_13924_ _26817_/Q _13919_/X _13912_/X _13923_/Y vssd1 vssd1 vccd1 vccd1 _26817_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17692_ _27413_/Q vssd1 vssd1 vccd1 vccd1 _17692_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19431_ _19431_/A vssd1 vssd1 vccd1 vccd1 _19431_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16643_ _16583_/A _16831_/B _16621_/A vssd1 vssd1 vccd1 vccd1 _16643_/X sky130_fd_sc_hd__o21ba_1
X_13855_ _13940_/B vssd1 vssd1 vccd1 vccd1 _13855_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19362_ _19362_/A _19362_/B _19362_/C vssd1 vssd1 vccd1 vccd1 _19363_/A sky130_fd_sc_hd__and3_1
X_16574_ _27403_/Q _16094_/X _16501_/X _14724_/A vssd1 vssd1 vccd1 vccd1 _16574_/X
+ sky130_fd_sc_hd__a22o_1
X_13786_ _26866_/Q _13778_/X _13780_/X _13785_/Y vssd1 vssd1 vccd1 vccd1 _26866_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18313_ _26957_/Q _26925_/Q _26893_/Q _26861_/Q _18244_/X _18269_/X vssd1 vssd1 vccd1
+ vccd1 _18313_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15525_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15534_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19293_ _19293_/A vssd1 vssd1 vccd1 vccd1 _26060_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18403_/A vssd1 vssd1 vccd1 vccd1 _18244_/X sky130_fd_sc_hd__buf_2
XFILLER_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15456_ _26244_/Q _13389_/X _15462_/S vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14407_ _26653_/Q _14405_/X _14398_/X _14406_/Y vssd1 vssd1 vccd1 vccd1 _26653_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18175_ _18358_/A vssd1 vssd1 vccd1 vccd1 _18175_/X sky130_fd_sc_hd__buf_2
XFILLER_117_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15387_ _15387_/A vssd1 vssd1 vccd1 vccd1 _26275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17126_ _17386_/S vssd1 vssd1 vccd1 vccd1 _17174_/S sky130_fd_sc_hd__clkbuf_2
X_14338_ _14344_/A vssd1 vssd1 vccd1 vccd1 _14393_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17057_ _17181_/A vssd1 vssd1 vccd1 vccd1 _17057_/X sky130_fd_sc_hd__clkbuf_2
X_14269_ _26704_/Q _14256_/X _14258_/X _14268_/Y vssd1 vssd1 vccd1 vccd1 _26704_/D
+ sky130_fd_sc_hd__a31o_1
X_16008_ _16136_/A vssd1 vssd1 vccd1 vccd1 _16132_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater301 _27649_/CLK vssd1 vssd1 vccd1 vccd1 _27654_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater312 _27705_/CLK vssd1 vssd1 vccd1 vccd1 _27706_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater323 _27770_/CLK vssd1 vssd1 vccd1 vccd1 _27711_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17959_ _17959_/A vssd1 vssd1 vccd1 vccd1 _17959_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater334 _27760_/CLK vssd1 vssd1 vccd1 vccd1 _27772_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater345 _27578_/CLK vssd1 vssd1 vccd1 vccd1 _27642_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_443 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater356 _27573_/CLK vssd1 vssd1 vccd1 vccd1 _27575_/CLK sky130_fd_sc_hd__clkbuf_1
X_20970_ _20970_/A vssd1 vssd1 vccd1 vccd1 _20970_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater367 _27682_/CLK vssd1 vssd1 vccd1 vccd1 _27411_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater378 _27559_/CLK vssd1 vssd1 vccd1 vccd1 _27452_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater389 _27196_/CLK vssd1 vssd1 vccd1 vccd1 _27462_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19629_ _19621_/X _19622_/X _19623_/X _19624_/X _19625_/X _19626_/X vssd1 vssd1 vccd1
+ vccd1 _19630_/A sky130_fd_sc_hd__mux4_1
XFILLER_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22640_ _22640_/A vssd1 vssd1 vccd1 vccd1 _22640_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22571_ _22561_/X _22562_/X _22563_/X _22564_/X _22565_/X _22566_/X vssd1 vssd1 vccd1
+ vccd1 _22572_/A sky130_fd_sc_hd__mux4_1
XFILLER_16_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21522_ _21522_/A vssd1 vssd1 vccd1 vccd1 _21522_/X sky130_fd_sc_hd__clkbuf_1
X_24310_ _16026_/X _16029_/Y _16033_/X _24217_/A vssd1 vssd1 vccd1 vccd1 _27439_/D
+ sky130_fd_sc_hd__a31oi_2
XFILLER_90_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25290_ _25299_/A _25290_/B vssd1 vssd1 vccd1 vccd1 _25291_/B sky130_fd_sc_hd__xnor2_1
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24241_ _24241_/A vssd1 vssd1 vccd1 vccd1 _27391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21453_ _21443_/X _21444_/X _21445_/X _21446_/X _21447_/X _21448_/X vssd1 vssd1 vccd1
+ vccd1 _21454_/A sky130_fd_sc_hd__mux4_1
XFILLER_147_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20404_ _20392_/X _20393_/X _20394_/X _20395_/X _20396_/X _20397_/X vssd1 vssd1 vccd1
+ vccd1 _20405_/A sky130_fd_sc_hd__mux4_1
X_24172_ _24172_/A vssd1 vssd1 vccd1 vccd1 _27357_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_21384_ _21384_/A vssd1 vssd1 vccd1 vccd1 _21384_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23123_ _23180_/S vssd1 vssd1 vccd1 vccd1 _23132_/S sky130_fd_sc_hd__clkbuf_2
X_20335_ _20335_/A vssd1 vssd1 vccd1 vccd1 _20335_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27931_ _27931_/A _15954_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
X_23054_ _23054_/A vssd1 vssd1 vccd1 vccd1 _27072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20266_ _20266_/A vssd1 vssd1 vccd1 vccd1 _20334_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22005_ _21997_/X _21998_/X _21999_/X _22000_/X _22002_/X _22004_/X vssd1 vssd1 vccd1
+ vccd1 _22006_/A sky130_fd_sc_hd__mux4_1
XFILLER_115_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20197_ _20197_/A vssd1 vssd1 vccd1 vccd1 _20197_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26813_ _22154_/X _26813_/D vssd1 vssd1 vccd1 vccd1 _26813_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27793_ _25628_/X _27793_/D vssd1 vssd1 vccd1 vccd1 _27793_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26744_ _21910_/X _26744_/D vssd1 vssd1 vccd1 vccd1 _26744_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23956_ _24003_/A vssd1 vssd1 vccd1 vccd1 _23956_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22907_ _22955_/A vssd1 vssd1 vccd1 vccd1 _22907_/X sky130_fd_sc_hd__clkbuf_1
X_26675_ _21680_/X _26675_/D vssd1 vssd1 vccd1 vccd1 _26675_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23887_ _27079_/Q _23860_/X _23861_/X _27111_/Q _23862_/X vssd1 vssd1 vccd1 vccd1
+ _23887_/X sky130_fd_sc_hd__a221o_1
XFILLER_44_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13640_ _13910_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13640_/Y sky130_fd_sc_hd__nor2_1
X_25626_ _25626_/A vssd1 vssd1 vccd1 vccd1 _27792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22838_ _22870_/A vssd1 vssd1 vccd1 vccd1 _22838_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25557_ _25592_/A vssd1 vssd1 vccd1 vccd1 _25557_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _27337_/Q _13022_/X _13030_/X _27305_/Q _13225_/X vssd1 vssd1 vccd1 vccd1
+ _14524_/A sky130_fd_sc_hd__a221oi_4
X_22769_ _22785_/A vssd1 vssd1 vccd1 vccd1 _22769_/X sky130_fd_sc_hd__clkbuf_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15310_ _15310_/A vssd1 vssd1 vccd1 vccd1 _26309_/D sky130_fd_sc_hd__clkbuf_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24508_ _24508_/A vssd1 vssd1 vccd1 vccd1 _27524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16287_/X _16288_/Y _16289_/X _16109_/A vssd1 vssd1 vccd1 vccd1 _16623_/B
+ sky130_fd_sc_hd__a31o_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25488_ _25487_/X _25461_/X _25462_/X _24863_/B _25463_/X vssd1 vssd1 vccd1 vccd1
+ _25488_/X sky130_fd_sc_hd__o311a_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27227_ _27302_/CLK _27227_/D vssd1 vssd1 vccd1 vccd1 _27227_/Q sky130_fd_sc_hd__dfxtp_1
X_15241_ _14782_/X _26339_/Q _15245_/S vssd1 vssd1 vccd1 vccd1 _15242_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24439_ _27618_/Q _24445_/B vssd1 vssd1 vccd1 vccd1 _24440_/A sky130_fd_sc_hd__and2_1
XFILLER_123_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27158_ _27852_/CLK _27158_/D vssd1 vssd1 vccd1 vccd1 _27158_/Q sky130_fd_sc_hd__dfxtp_1
X_15172_ _15172_/A vssd1 vssd1 vccd1 vccd1 _26370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14123_ _14388_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26109_ _19693_/X _26109_/D vssd1 vssd1 vccd1 vccd1 _26109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19980_ _19972_/X _19973_/X _19974_/X _19975_/X _19976_/X _19977_/X vssd1 vssd1 vccd1
+ vccd1 _19981_/A sky130_fd_sc_hd__mux4_1
X_27089_ _27121_/CLK _27089_/D vssd1 vssd1 vccd1 vccd1 _27089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18931_ _26269_/Q _26237_/Q _26205_/Q _26173_/Q _18778_/X _18930_/X vssd1 vssd1 vccd1
+ vccd1 _18931_/X sky130_fd_sc_hd__mux4_2
XFILLER_107_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14054_ _26780_/Q _14042_/X _14038_/X _14053_/Y vssd1 vssd1 vccd1 vccd1 _26780_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _27796_/Q _13009_/B vssd1 vssd1 vccd1 vccd1 _13006_/A sky130_fd_sc_hd__and2_1
X_18862_ _26395_/Q _26363_/Q _26331_/Q _26299_/Q _18824_/X _18826_/X vssd1 vssd1 vccd1
+ vccd1 _18862_/X sky130_fd_sc_hd__mux4_1
X_17813_ _18156_/A vssd1 vssd1 vccd1 vccd1 _17813_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18793_ _19465_/A vssd1 vssd1 vccd1 vccd1 _18793_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17744_ _27429_/Q vssd1 vssd1 vccd1 vccd1 _17744_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14956_ _14956_/A vssd1 vssd1 vccd1 vccd1 _26458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13907_ _13920_/A vssd1 vssd1 vccd1 vccd1 _13917_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17675_ _18691_/A _23182_/B _23109_/A vssd1 vssd1 vccd1 vccd1 _17757_/A sky130_fd_sc_hd__and3b_2
X_14887_ _14955_/S vssd1 vssd1 vccd1 vccd1 _14896_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_165_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19414_ _19414_/A vssd1 vssd1 vccd1 vccd1 _19414_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16626_ _16626_/A vssd1 vssd1 vccd1 vccd1 _16626_/X sky130_fd_sc_hd__clkbuf_2
X_13838_ _13930_/A _13838_/B vssd1 vssd1 vccd1 vccd1 _13838_/Y sky130_fd_sc_hd__nor2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19345_ _27814_/Q _26575_/Q _26447_/Q _26127_/Q _19255_/X _19321_/X vssd1 vssd1 vccd1
+ vccd1 _19345_/X sky130_fd_sc_hd__mux4_2
XFILLER_189_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16557_ _27401_/Q _16557_/B vssd1 vssd1 vccd1 vccd1 _16557_/Y sky130_fd_sc_hd__nand2_1
X_13769_ _26872_/Q _13761_/X _13764_/X _13768_/Y vssd1 vssd1 vccd1 vccd1 _26872_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _13128_/X _26221_/Q _15512_/S vssd1 vssd1 vccd1 vccd1 _15509_/A sky130_fd_sc_hd__mux2_1
X_19276_ _26956_/Q _26924_/Q _26892_/Q _26860_/Q _19208_/X _19253_/X vssd1 vssd1 vccd1
+ vccd1 _19276_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16488_ _16497_/B _16489_/C _16670_/A vssd1 vssd1 vccd1 vccd1 _16493_/B sky130_fd_sc_hd__a21o_1
XFILLER_148_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18227_ _17995_/X _18222_/X _18224_/X _18226_/X _18016_/X vssd1 vssd1 vccd1 vccd1
+ _18240_/B sky130_fd_sc_hd__a221o_1
X_15439_ _15439_/A vssd1 vssd1 vccd1 vccd1 _26252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_702 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18158_ _18057_/X _18154_/X _18157_/X _18062_/X vssd1 vssd1 vccd1 vccd1 _18158_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17109_ _25819_/Q _26018_/Q _17158_/S vssd1 vssd1 vccd1 vccd1 _17109_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18089_ _26531_/Q _26499_/Q _26467_/Q _27043_/Q _17899_/X _17901_/X vssd1 vssd1 vccd1
+ vccd1 _18089_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20120_ _20114_/X _20115_/X _20116_/X _20117_/X _20118_/X _20119_/X vssd1 vssd1 vccd1
+ vccd1 _20121_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20051_ _20051_/A vssd1 vssd1 vccd1 vccd1 _20051_/X sky130_fd_sc_hd__clkbuf_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater120 _27675_/CLK vssd1 vssd1 vccd1 vccd1 _27678_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater131 _27094_/CLK vssd1 vssd1 vccd1 vccd1 _26039_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater142 _27127_/CLK vssd1 vssd1 vccd1 vccd1 _27115_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23810_ _24047_/S vssd1 vssd1 vccd1 vccd1 _23846_/S sky130_fd_sc_hd__clkbuf_2
Xrepeater153 _27789_/CLK vssd1 vssd1 vccd1 vccd1 _27418_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24790_ _24790_/A _24800_/B vssd1 vssd1 vccd1 vccd1 _24790_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater164 _27130_/CLK vssd1 vssd1 vccd1 vccd1 _27827_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater175 _27077_/CLK vssd1 vssd1 vccd1 vccd1 _26022_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater186 _27416_/CLK vssd1 vssd1 vccd1 vccd1 _27414_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _14507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23741_ _27785_/Q vssd1 vssd1 vccd1 vccd1 _23777_/A sky130_fd_sc_hd__clkbuf_2
X_20953_ _20953_/A vssd1 vssd1 vccd1 vccd1 _20953_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater197 _26012_/CLK vssd1 vssd1 vccd1 vccd1 _27676_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26460_ _20928_/X _26460_/D vssd1 vssd1 vccd1 vccd1 _26460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _20884_/A vssd1 vssd1 vccd1 vccd1 _20884_/X sky130_fd_sc_hd__clkbuf_1
X_23672_ _24862_/A _27242_/Q _23672_/S vssd1 vssd1 vccd1 vccd1 _23673_/A sky130_fd_sc_hd__mux2_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25411_ _27744_/Q input56/X _25413_/S vssd1 vssd1 vccd1 vccd1 _25412_/A sky130_fd_sc_hd__mux2_1
X_22623_ _22609_/X _22610_/X _22611_/X _22612_/X _22615_/X _22618_/X vssd1 vssd1 vccd1
+ vccd1 _22624_/A sky130_fd_sc_hd__mux4_1
X_26391_ _20677_/X _26391_/D vssd1 vssd1 vccd1 vccd1 _26391_/Q sky130_fd_sc_hd__dfxtp_1
X_22554_ _22554_/A vssd1 vssd1 vccd1 vccd1 _22554_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25342_ _25342_/A _25341_/Y vssd1 vssd1 vccd1 vccd1 _25343_/B sky130_fd_sc_hd__or2b_1
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21505_ _21494_/X _21496_/X _21498_/X _21500_/X _21501_/X _21502_/X vssd1 vssd1 vccd1
+ vccd1 _21506_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22485_ _22471_/X _22472_/X _22473_/X _22474_/X _22475_/X _22476_/X vssd1 vssd1 vccd1
+ vccd1 _22486_/A sky130_fd_sc_hd__mux4_1
X_25273_ _25273_/A _25273_/B vssd1 vssd1 vccd1 vccd1 _25274_/B sky130_fd_sc_hd__or2_1
X_27012_ _22848_/X _27012_/D vssd1 vssd1 vccd1 vccd1 _27012_/Q sky130_fd_sc_hd__dfxtp_1
X_21436_ _21436_/A vssd1 vssd1 vccd1 vccd1 _21436_/X sky130_fd_sc_hd__clkbuf_1
X_24224_ _24304_/A vssd1 vssd1 vccd1 vccd1 _24235_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24155_ _24155_/A vssd1 vssd1 vccd1 vccd1 _27349_/D sky130_fd_sc_hd__clkbuf_1
X_21367_ _21357_/X _21358_/X _21359_/X _21360_/X _21361_/X _21362_/X vssd1 vssd1 vccd1
+ vccd1 _21368_/A sky130_fd_sc_hd__mux4_1
XFILLER_123_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23106_ _23106_/A vssd1 vssd1 vccd1 vccd1 _27096_/D sky130_fd_sc_hd__clkbuf_1
X_20318_ _20334_/A vssd1 vssd1 vccd1 vccd1 _20318_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24086_ _24119_/A vssd1 vssd1 vccd1 vccd1 _24095_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_21298_ _21298_/A vssd1 vssd1 vccd1 vccd1 _21298_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23037_ _27375_/Q _24001_/A vssd1 vssd1 vccd1 vccd1 _23094_/A sky130_fd_sc_hd__and2_1
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20249_ _20249_/A vssd1 vssd1 vccd1 vccd1 _20249_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27845_ _27845_/CLK _27845_/D vssd1 vssd1 vccd1 vccd1 _27845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14810_ _14810_/A vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27776_ _27776_/CLK _27776_/D vssd1 vssd1 vccd1 vccd1 _27776_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15790_ _13067_/X _26103_/Q _15794_/S vssd1 vssd1 vccd1 vccd1 _15791_/A sky130_fd_sc_hd__mux2_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24988_ _25075_/A vssd1 vssd1 vccd1 vccd1 _25024_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_92_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26727_ _21858_/X _26727_/D vssd1 vssd1 vccd1 vccd1 _26727_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14741_ _14740_/X _26544_/Q _14741_/S vssd1 vssd1 vccd1 vccd1 _14742_/A sky130_fd_sc_hd__mux2_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23939_ _27085_/Q _27117_/Q _23939_/S vssd1 vssd1 vccd1 vccd1 _23939_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _27419_/Q vssd1 vssd1 vccd1 vccd1 _17460_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26658_ _21612_/X _26658_/D vssd1 vssd1 vccd1 vccd1 _26658_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _15745_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14672_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16411_ _16711_/A _16411_/B vssd1 vssd1 vccd1 vccd1 _16710_/A sky130_fd_sc_hd__xnor2_1
X_13623_ _13649_/A vssd1 vssd1 vccd1 vccd1 _13634_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25609_ _27719_/Q _25433_/X _25435_/X vssd1 vssd1 vccd1 vccd1 _25609_/Y sky130_fd_sc_hd__a21oi_1
X_17391_ _25653_/A vssd1 vssd1 vccd1 vccd1 _19830_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_26589_ _21372_/X _26589_/D vssd1 vssd1 vccd1 vccd1 _26589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19130_ _19222_/A _19130_/B _19130_/C vssd1 vssd1 vccd1 vccd1 _19131_/A sky130_fd_sc_hd__and3_1
XFILLER_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16342_ _16342_/A _16353_/A vssd1 vssd1 vccd1 vccd1 _16342_/Y sky130_fd_sc_hd__nor2_1
XFILLER_198_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _27341_/Q _13529_/X _13530_/X _27309_/Q _13201_/X vssd1 vssd1 vccd1 vccd1
+ _14511_/A sky130_fd_sc_hd__a221oi_4
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_753 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater78 _27430_/CLK vssd1 vssd1 vccd1 vccd1 _27151_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater89 _27849_/CLK vssd1 vssd1 vccd1 vccd1 _27153_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_146_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19061_ _19401_/A vssd1 vssd1 vccd1 vccd1 _19061_/X sky130_fd_sc_hd__clkbuf_4
X_16273_ _16108_/A _16268_/X _16270_/Y _16271_/X _16272_/X vssd1 vssd1 vccd1 vccd1
+ _16809_/A sky130_fd_sc_hd__o41a_1
XFILLER_173_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13485_ _13887_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13485_/Y sky130_fd_sc_hd__nor2_1
XFILLER_201_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1021 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18012_ _18012_/A vssd1 vssd1 vccd1 vccd1 _24388_/A sky130_fd_sc_hd__buf_4
X_15224_ _15224_/A vssd1 vssd1 vccd1 vccd1 _26347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15155_ _15155_/A vssd1 vssd1 vccd1 vccd1 _26378_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ _26763_/Q _14104_/X _14093_/X _14105_/Y vssd1 vssd1 vccd1 vccd1 _26763_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_181_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19963_ _19963_/A vssd1 vssd1 vccd1 vccd1 _19963_/X sky130_fd_sc_hd__clkbuf_1
X_15086_ _14766_/X _26408_/Q _15090_/S vssd1 vssd1 vccd1 vccd1 _15087_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14037_ _26785_/Q _14024_/X _14019_/X _14036_/Y vssd1 vssd1 vccd1 vccd1 _26785_/D
+ sky130_fd_sc_hd__a31o_1
X_18914_ _19165_/A vssd1 vssd1 vccd1 vccd1 _18930_/A sky130_fd_sc_hd__buf_4
XFILLER_171_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19894_ _19882_/X _19883_/X _19884_/X _19885_/X _19886_/X _19887_/X vssd1 vssd1 vccd1
+ vccd1 _19895_/A sky130_fd_sc_hd__mux4_1
XFILLER_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18845_ _26811_/Q _26779_/Q _26747_/Q _26715_/Q _18767_/X _18770_/X vssd1 vssd1 vccd1
+ vccd1 _18846_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18776_ _18828_/A vssd1 vssd1 vccd1 vccd1 _18922_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15988_ _15988_/A vssd1 vssd1 vccd1 vccd1 _15988_/Y sky130_fd_sc_hd__inv_2
X_17727_ _17727_/A vssd1 vssd1 vccd1 vccd1 _25927_/D sky130_fd_sc_hd__clkbuf_1
X_14939_ _14939_/A vssd1 vssd1 vccd1 vccd1 _26466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17658_ _17658_/A vssd1 vssd1 vccd1 vccd1 _17667_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_51_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16609_ _16609_/A _16609_/B vssd1 vssd1 vccd1 vccd1 _16610_/B sky130_fd_sc_hd__nand2_1
X_17589_ _17508_/X _25869_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17590_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19328_ _19419_/A _19328_/B vssd1 vssd1 vccd1 vccd1 _19328_/X sky130_fd_sc_hd__or2_1
XFILLER_91_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19259_ _19250_/X _19252_/X _19257_/X _19186_/X _19258_/X vssd1 vssd1 vccd1 vccd1
+ _19268_/B sky130_fd_sc_hd__a221o_1
XFILLER_137_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22270_ _22270_/A vssd1 vssd1 vccd1 vccd1 _22270_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21221_ _21211_/X _21212_/X _21213_/X _21214_/X _21216_/X _21218_/X vssd1 vssd1 vccd1
+ vccd1 _21222_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21152_ _21200_/A vssd1 vssd1 vccd1 vccd1 _21152_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20103_ _20151_/A vssd1 vssd1 vccd1 vccd1 _20103_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25960_ _25969_/CLK _25960_/D vssd1 vssd1 vccd1 vccd1 _25960_/Q sky130_fd_sc_hd__dfxtp_1
X_21083_ _21077_/X _21078_/X _21079_/X _21080_/X _21081_/X _21082_/X vssd1 vssd1 vccd1
+ vccd1 _21084_/A sky130_fd_sc_hd__mux4_1
XFILLER_59_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24911_ _24906_/A _24910_/C _27772_/Q vssd1 vssd1 vccd1 vccd1 _24912_/B sky130_fd_sc_hd__a21oi_1
X_20034_ _20028_/X _20029_/X _20030_/X _20031_/X _20032_/X _20033_/X vssd1 vssd1 vccd1
+ vccd1 _20035_/A sky130_fd_sc_hd__mux4_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25891_ _27842_/CLK _25891_/D vssd1 vssd1 vccd1 vccd1 _25891_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27630_ _27633_/CLK _27630_/D vssd1 vssd1 vccd1 vccd1 _27630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24842_ _24935_/A vssd1 vssd1 vccd1 vccd1 _24863_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27561_ _27562_/CLK _27561_/D vssd1 vssd1 vccd1 vccd1 _27561_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24773_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24773_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21985_ _21985_/A vssd1 vssd1 vccd1 vccd1 _21985_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26512_ _21104_/X _26512_/D vssd1 vssd1 vccd1 vccd1 _26512_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23724_ _24063_/A vssd1 vssd1 vccd1 vccd1 _24005_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27492_ _27612_/CLK _27492_/D vssd1 vssd1 vccd1 vccd1 _27492_/Q sky130_fd_sc_hd__dfxtp_1
X_20936_ _20936_/A vssd1 vssd1 vccd1 vccd1 _20936_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26443_ _20861_/X _26443_/D vssd1 vssd1 vccd1 vccd1 _26443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20867_ _20867_/A vssd1 vssd1 vccd1 vccd1 _20867_/X sky130_fd_sc_hd__clkbuf_1
X_23655_ _25977_/Q _27234_/Q _23661_/S vssd1 vssd1 vccd1 vccd1 _23656_/A sky130_fd_sc_hd__mux2_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22606_ _22606_/A vssd1 vssd1 vccd1 vccd1 _22606_/X sky130_fd_sc_hd__clkbuf_1
X_26374_ _20615_/X _26374_/D vssd1 vssd1 vccd1 vccd1 _26374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23586_ _23596_/A _23586_/B vssd1 vssd1 vccd1 vccd1 _23587_/A sky130_fd_sc_hd__and2_1
XFILLER_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20798_ _21147_/A vssd1 vssd1 vccd1 vccd1 _20866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_168_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25325_ _25325_/A _25325_/B vssd1 vssd1 vccd1 vccd1 _25326_/B sky130_fd_sc_hd__xnor2_1
XFILLER_168_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22537_ _22537_/A vssd1 vssd1 vccd1 vccd1 _22887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_195_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28001__467 vssd1 vssd1 vccd1 vccd1 _28001__467/HI _28001_/A sky130_fd_sc_hd__conb_1
X_25256_ _27538_/Q _27506_/Q vssd1 vssd1 vccd1 vccd1 _25267_/B sky130_fd_sc_hd__nor2_1
X_13270_ _13270_/A vssd1 vssd1 vccd1 vccd1 _27024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22468_ _22468_/A vssd1 vssd1 vccd1 vccd1 _22468_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24207_ _24207_/A _24210_/B vssd1 vssd1 vccd1 vccd1 _27371_/D sky130_fd_sc_hd__nor2_1
X_21419_ _21408_/X _21410_/X _21412_/X _21414_/X _21415_/X _21416_/X vssd1 vssd1 vccd1
+ vccd1 _21420_/A sky130_fd_sc_hd__mux4_1
XFILLER_5_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22399_ _22385_/X _22386_/X _22387_/X _22388_/X _22389_/X _22390_/X vssd1 vssd1 vccd1
+ vccd1 _22400_/A sky130_fd_sc_hd__mux4_1
X_25187_ _27529_/Q _27497_/Q vssd1 vssd1 vccd1 vccd1 _25187_/X sky130_fd_sc_hd__or2_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24138_ _27447_/Q _24140_/B vssd1 vssd1 vccd1 vccd1 _24139_/A sky130_fd_sc_hd__and2_1
XFILLER_155_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16960_ _16960_/A vssd1 vssd1 vccd1 vccd1 _16982_/C sky130_fd_sc_hd__clkbuf_1
X_24069_ _24069_/A vssd1 vssd1 vccd1 vccd1 _27311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _15912_/A vssd1 vssd1 vccd1 vccd1 _15911_/Y sky130_fd_sc_hd__inv_2
X_16891_ _16890_/A _16890_/C _16890_/B vssd1 vssd1 vccd1 vccd1 _16891_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18630_ _25982_/Q _17689_/X _18630_/S vssd1 vssd1 vccd1 vccd1 _18631_/A sky130_fd_sc_hd__mux2_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15842_ _15842_/A vssd1 vssd1 vccd1 vccd1 _26080_/D sky130_fd_sc_hd__clkbuf_1
X_27828_ _27830_/CLK _27828_/D vssd1 vssd1 vccd1 vccd1 _27828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18561_ _26424_/Q _26392_/Q _26360_/Q _26328_/Q _18462_/X _18486_/X vssd1 vssd1 vccd1
+ vccd1 _18561_/X sky130_fd_sc_hd__mux4_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15773_/A vssd1 vssd1 vccd1 vccd1 _23562_/A sky130_fd_sc_hd__clkbuf_4
X_27759_ _27760_/CLK _27759_/D vssd1 vssd1 vccd1 vccd1 _27759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ _27805_/Q _12987_/B vssd1 vssd1 vccd1 vccd1 _12986_/A sky130_fd_sc_hd__and2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17512_ _17511_/X _25838_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__mux2_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _14724_/A vssd1 vssd1 vccd1 vccd1 _14724_/X sky130_fd_sc_hd__clkbuf_4
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _18492_/A vssd1 vssd1 vccd1 vccd1 _25970_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17443_ _17443_/A vssd1 vssd1 vccd1 vccd1 _25816_/D sky130_fd_sc_hd__clkbuf_1
X_14655_ _26575_/Q _14645_/X _14653_/X _14654_/Y vssd1 vssd1 vccd1 vccd1 _26575_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _13876_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13606_/Y sky130_fd_sc_hd__nor2_1
X_17374_ _17116_/A _17369_/X _17371_/X _17373_/X vssd1 vssd1 vccd1 vccd1 _17374_/X
+ sky130_fd_sc_hd__o22a_1
X_14586_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14597_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19113_ _19113_/A _19113_/B vssd1 vssd1 vccd1 vccd1 _19113_/X sky130_fd_sc_hd__or2_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16325_ _16752_/B vssd1 vssd1 vccd1 vccd1 _16754_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13537_ _14497_/A vssd1 vssd1 vccd1 vccd1 _13915_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19044_ _19208_/A vssd1 vssd1 vccd1 vccd1 _19044_/X sky130_fd_sc_hd__clkbuf_4
X_16256_ _16422_/A _16256_/B _16256_/C _16255_/Y vssd1 vssd1 vccd1 vccd1 _16257_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_139_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13468_ _26963_/Q _13464_/X _13457_/X _13467_/Y vssd1 vssd1 vccd1 vccd1 _26963_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15207_ _15207_/A vssd1 vssd1 vccd1 vccd1 _26355_/D sky130_fd_sc_hd__clkbuf_1
X_16187_ _16180_/X _16182_/X _16185_/X _16186_/X vssd1 vssd1 vccd1 vccd1 _16200_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13399_ _26977_/Q _13398_/X _13399_/S vssd1 vssd1 vccd1 vccd1 _13400_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _26385_/Q _13347_/X _15140_/S vssd1 vssd1 vccd1 vccd1 _15139_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19946_ _19940_/X _19941_/X _19942_/X _19943_/X _19944_/X _19945_/X vssd1 vssd1 vccd1
+ vccd1 _19947_/A sky130_fd_sc_hd__mux4_1
X_15069_ _15069_/A vssd1 vssd1 vccd1 vccd1 _26416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19877_ _19877_/A vssd1 vssd1 vccd1 vccd1 _19877_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18828_ _18828_/A vssd1 vssd1 vccd1 vccd1 _19414_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18759_ _26040_/Q _17772_/X _18761_/S vssd1 vssd1 vccd1 vccd1 _18760_/A sky130_fd_sc_hd__mux2_1
X_21770_ _21770_/A vssd1 vssd1 vccd1 vccd1 _21770_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20721_ _20721_/A vssd1 vssd1 vccd1 vccd1 _20721_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20652_ _20684_/A vssd1 vssd1 vccd1 vccd1 _20652_/X sky130_fd_sc_hd__clkbuf_1
X_23440_ _27170_/Q _23443_/B vssd1 vssd1 vccd1 vccd1 _23440_/X sky130_fd_sc_hd__or2_1
XFILLER_196_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23371_ _27771_/Q vssd1 vssd1 vccd1 vccd1 _24780_/A sky130_fd_sc_hd__inv_2
X_20583_ _20599_/A vssd1 vssd1 vccd1 vccd1 _20583_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25110_ _25733_/A _25110_/B vssd1 vssd1 vccd1 vccd1 _25143_/A sky130_fd_sc_hd__nand2_1
X_22322_ _22322_/A vssd1 vssd1 vccd1 vccd1 _22322_/X sky130_fd_sc_hd__clkbuf_1
X_26090_ _19628_/X _26090_/D vssd1 vssd1 vccd1 vccd1 _26090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22253_ _22245_/X _22246_/X _22247_/X _22248_/X _22249_/X _22250_/X vssd1 vssd1 vccd1
+ vccd1 _22254_/A sky130_fd_sc_hd__mux4_1
X_25041_ _25038_/X _25039_/X _25074_/S vssd1 vssd1 vccd1 vccd1 _25041_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21204_ _21204_/A vssd1 vssd1 vccd1 vccd1 _21204_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22184_ _22184_/A vssd1 vssd1 vccd1 vccd1 _22184_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_535 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21135_ _21125_/X _21126_/X _21127_/X _21128_/X _21130_/X _21132_/X vssd1 vssd1 vccd1
+ vccd1 _21136_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26992_ _22778_/X _26992_/D vssd1 vssd1 vccd1 vccd1 _26992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25943_ _27110_/CLK _25943_/D vssd1 vssd1 vccd1 vccd1 _25943_/Q sky130_fd_sc_hd__dfxtp_1
X_21066_ _21114_/A vssd1 vssd1 vccd1 vccd1 _21066_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20017_ _20065_/A vssd1 vssd1 vccd1 vccd1 _20017_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25874_ _27857_/CLK _25874_/D vssd1 vssd1 vccd1 vccd1 _25874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27613_ _27614_/CLK _27613_/D vssd1 vssd1 vccd1 vccd1 _27613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24825_ _24825_/A _25601_/B vssd1 vssd1 vccd1 vccd1 _24825_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27544_ _27667_/CLK _27544_/D vssd1 vssd1 vccd1 vccd1 _27544_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24756_ _24756_/A _24759_/B vssd1 vssd1 vccd1 vccd1 _24756_/Y sky130_fd_sc_hd__nand2_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ _22000_/A vssd1 vssd1 vccd1 vccd1 _21968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23707_ _23707_/A vssd1 vssd1 vccd1 vccd1 _23716_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27475_ _27475_/CLK _27475_/D vssd1 vssd1 vccd1 vccd1 _27475_/Q sky130_fd_sc_hd__dfxtp_1
X_20919_ _20905_/X _20906_/X _20907_/X _20908_/X _20909_/X _20910_/X vssd1 vssd1 vccd1
+ vccd1 _20920_/A sky130_fd_sc_hd__mux4_1
X_24687_ _24700_/A vssd1 vssd1 vccd1 vccd1 _24687_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _21899_/A vssd1 vssd1 vccd1 vccd1 _21899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14440_ _26644_/Q _14421_/X _14437_/X _14439_/Y vssd1 vssd1 vccd1 vccd1 _26644_/D
+ sky130_fd_sc_hd__a31o_1
X_26426_ _20809_/X _26426_/D vssd1 vssd1 vccd1 vccd1 _26426_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23638_ _23638_/A _23638_/B _23638_/C vssd1 vssd1 vccd1 vccd1 _23638_/X sky130_fd_sc_hd__and3_1
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _14398_/A vssd1 vssd1 vccd1 vccd1 _14371_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26357_ _20561_/X _26357_/D vssd1 vssd1 vccd1 vccd1 _26357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23569_ _23569_/A vssd1 vssd1 vccd1 vccd1 _27211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16110_ _16110_/A vssd1 vssd1 vccd1 vccd1 _16151_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25308_ _25308_/A vssd1 vssd1 vccd1 vccd1 _25308_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _13421_/S vssd1 vssd1 vccd1 vccd1 _13335_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17090_ _17088_/X _17089_/X _17113_/S vssd1 vssd1 vccd1 vccd1 _17090_/X sky130_fd_sc_hd__mux2_1
X_26288_ _20315_/X _26288_/D vssd1 vssd1 vccd1 vccd1 _26288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16041_ _27474_/Q _27370_/Q vssd1 vssd1 vccd1 vccd1 _16041_/X sky130_fd_sc_hd__or2b_1
X_25239_ _27536_/Q _27504_/Q vssd1 vssd1 vccd1 vccd1 _25241_/A sky130_fd_sc_hd__nand2_1
X_13253_ _13253_/A vssd1 vssd1 vccd1 vccd1 _27032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13184_ _16235_/A vssd1 vssd1 vccd1 vccd1 _13184_/X sky130_fd_sc_hd__buf_2
XFILLER_124_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19800_ _19800_/A vssd1 vssd1 vccd1 vccd1 _19800_/X sky130_fd_sc_hd__clkbuf_2
X_17992_ _18028_/A _17992_/B _17992_/C vssd1 vssd1 vccd1 vccd1 _17993_/A sky130_fd_sc_hd__and3_1
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19731_ _19800_/A vssd1 vssd1 vccd1 vccd1 _19731_/X sky130_fd_sc_hd__clkbuf_2
X_16943_ _19448_/A _27487_/Q _27486_/Q _18945_/A _16942_/X vssd1 vssd1 vccd1 vccd1
+ _16943_/X sky130_fd_sc_hd__o221a_1
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16874_ _24242_/A _25618_/A _16874_/C _16874_/D vssd1 vssd1 vccd1 vccd1 _16875_/D
+ sky130_fd_sc_hd__and4_1
X_19662_ _19834_/A vssd1 vssd1 vccd1 vccd1 _19728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18613_ _18613_/A _18613_/B vssd1 vssd1 vccd1 vccd1 _25115_/A sky130_fd_sc_hd__xor2_1
X_15825_ _13161_/X _26087_/Q _15827_/S vssd1 vssd1 vccd1 vccd1 _15826_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19593_ _19625_/A vssd1 vssd1 vccd1 vccd1 _19593_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15756_/A _15758_/B vssd1 vssd1 vccd1 vccd1 _15756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18544_ _18542_/X _18543_/X _18580_/S vssd1 vssd1 vccd1 vccd1 _18544_/X sky130_fd_sc_hd__mux2_2
X_12968_ _27813_/Q _12976_/B vssd1 vssd1 vccd1 vccd1 _12969_/A sky130_fd_sc_hd__and2_1
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _15781_/A _14707_/B vssd1 vssd1 vccd1 vccd1 _14707_/Y sky130_fd_sc_hd__nor2_1
X_18475_ _18475_/A _18474_/X vssd1 vssd1 vccd1 vccd1 _18475_/X sky130_fd_sc_hd__or2b_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15687_ _13222_/X _26141_/Q _15689_/S vssd1 vssd1 vccd1 vccd1 _15688_/A sky130_fd_sc_hd__mux2_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_370 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_381 _13222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _17408_/X _25811_/Q _17438_/S vssd1 vssd1 vccd1 vccd1 _17427_/A sky130_fd_sc_hd__mux2_1
X_14638_ _26581_/Q _14630_/X _14624_/X _14637_/Y vssd1 vssd1 vccd1 vccd1 _26581_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17357_ _27223_/Q _17356_/X _17367_/S vssd1 vssd1 vccd1 vccd1 _17358_/A sky130_fd_sc_hd__mux2_1
X_14569_ _15730_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14569_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _16308_/A _16308_/B vssd1 vssd1 vccd1 vccd1 _16309_/B sky130_fd_sc_hd__or2_1
X_17288_ _27849_/Q _27153_/Q _25898_/Q _25866_/Q _17264_/X _17252_/X vssd1 vssd1 vccd1
+ vccd1 _17288_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19027_ _19123_/A _19027_/B vssd1 vssd1 vccd1 vccd1 _19027_/X sky130_fd_sc_hd__or2_1
X_16239_ _16428_/A _16358_/A _16407_/A _16447_/D vssd1 vssd1 vccd1 vccd1 _16256_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27993__459 vssd1 vssd1 vccd1 vccd1 _27993__459/HI _27993_/A sky130_fd_sc_hd__conb_1
XFILLER_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19929_ _19977_/A vssd1 vssd1 vccd1 vccd1 _19929_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22940_ _22956_/A vssd1 vssd1 vccd1 vccd1 _22940_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22871_ _22871_/A vssd1 vssd1 vccd1 vccd1 _22871_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24610_ _24610_/A vssd1 vssd1 vccd1 vccd1 _27564_/D sky130_fd_sc_hd__clkbuf_1
X_21822_ _21822_/A vssd1 vssd1 vccd1 vccd1 _21822_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25590_ _18594_/A _25321_/B _25589_/X _25566_/X vssd1 vssd1 vccd1 vccd1 _25590_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24541_ _24541_/A vssd1 vssd1 vccd1 vccd1 _27534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21753_ _21737_/X _21738_/X _21739_/X _21740_/X _21743_/X _21746_/X vssd1 vssd1 vccd1
+ vccd1 _21754_/A sky130_fd_sc_hd__mux4_1
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20704_ _20704_/A vssd1 vssd1 vccd1 vccd1 _20771_/A sky130_fd_sc_hd__buf_2
X_27260_ _27778_/CLK _27260_/D vssd1 vssd1 vccd1 vccd1 _27260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24472_ _27633_/Q _24478_/B vssd1 vssd1 vccd1 vccd1 _24473_/A sky130_fd_sc_hd__and2_1
X_21684_ _21684_/A vssd1 vssd1 vccd1 vccd1 _21684_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26211_ _20053_/X _26211_/D vssd1 vssd1 vccd1 vccd1 _26211_/Q sky130_fd_sc_hd__dfxtp_1
X_23423_ _27163_/Q _23430_/B vssd1 vssd1 vccd1 vccd1 _23423_/X sky130_fd_sc_hd__or2_1
X_20635_ _20635_/A vssd1 vssd1 vccd1 vccd1 _20635_/X sky130_fd_sc_hd__clkbuf_1
X_27191_ _27607_/CLK _27191_/D vssd1 vssd1 vccd1 vccd1 _27191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26142_ _19807_/X _26142_/D vssd1 vssd1 vccd1 vccd1 _26142_/Q sky130_fd_sc_hd__dfxtp_1
X_23354_ _27255_/Q vssd1 vssd1 vccd1 vccd1 _23354_/Y sky130_fd_sc_hd__inv_2
X_20566_ _20598_/A vssd1 vssd1 vccd1 vccd1 _20566_/X sky130_fd_sc_hd__clkbuf_1
X_22305_ _22299_/X _22300_/X _22301_/X _22302_/X _22303_/X _22304_/X vssd1 vssd1 vccd1
+ vccd1 _22306_/A sky130_fd_sc_hd__mux4_1
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26073_ _26073_/CLK _26073_/D vssd1 vssd1 vccd1 vccd1 _26073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23285_ input56/X vssd1 vssd1 vccd1 vccd1 _23285_/Y sky130_fd_sc_hd__inv_2
X_20497_ _20513_/A vssd1 vssd1 vccd1 vccd1 _20497_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25024_ _27968_/A _25023_/X _25024_/S vssd1 vssd1 vccd1 vccd1 _25025_/A sky130_fd_sc_hd__mux2_1
X_22236_ _22236_/A vssd1 vssd1 vccd1 vccd1 _22236_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22167_ _22157_/X _22158_/X _22159_/X _22160_/X _22161_/X _22162_/X vssd1 vssd1 vccd1
+ vccd1 _22168_/A sky130_fd_sc_hd__mux4_1
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21118_ _21118_/A vssd1 vssd1 vccd1 vccd1 _21118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22098_ _22098_/A vssd1 vssd1 vccd1 vccd1 _22098_/X sky130_fd_sc_hd__clkbuf_1
X_26975_ _22726_/X _26975_/D vssd1 vssd1 vccd1 vccd1 _26975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _13940_/A _13940_/B vssd1 vssd1 vccd1 vccd1 _13940_/Y sky130_fd_sc_hd__nor2_1
X_25926_ _25991_/CLK _25926_/D vssd1 vssd1 vccd1 vccd1 _25926_/Q sky130_fd_sc_hd__dfxtp_1
X_21049_ _21039_/X _21040_/X _21041_/X _21042_/X _21044_/X _21046_/X vssd1 vssd1 vccd1
+ vccd1 _21050_/A sky130_fd_sc_hd__mux4_1
XFILLER_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_474 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13871_ _26837_/Q _13865_/X _13855_/X _13870_/Y vssd1 vssd1 vccd1 vccd1 _26837_/D
+ sky130_fd_sc_hd__a31o_1
X_25857_ _27144_/CLK _25857_/D vssd1 vssd1 vccd1 vccd1 _25857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15610_ _15610_/A vssd1 vssd1 vccd1 vccd1 _26176_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1096 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24808_ _24808_/A _24815_/B vssd1 vssd1 vccd1 vccd1 _24808_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16590_ _27404_/Q _16312_/X _16501_/X _14721_/A vssd1 vssd1 vccd1 vccd1 _16590_/X
+ sky130_fd_sc_hd__a22o_1
X_25788_ _17498_/X _27849_/Q _25790_/S vssd1 vssd1 vccd1 vccd1 _25789_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27527_ _27527_/CLK _27527_/D vssd1 vssd1 vccd1 vccd1 _27527_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _13216_/X _26206_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15542_/A sky130_fd_sc_hd__mux2_1
X_24739_ _24835_/A vssd1 vssd1 vccd1 vccd1 _24740_/A sky130_fd_sc_hd__inv_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _26538_/Q _26506_/Q _26474_/Q _27050_/Q _18233_/X _18259_/X vssd1 vssd1 vccd1
+ vccd1 _18260_/X sky130_fd_sc_hd__mux4_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27458_ _27458_/CLK _27458_/D vssd1 vssd1 vccd1 vccd1 _27458_/Q sky130_fd_sc_hd__dfxtp_1
X_15472_ _15472_/A vssd1 vssd1 vccd1 vccd1 _26237_/D sky130_fd_sc_hd__clkbuf_1
X_28007__473 vssd1 vssd1 vccd1 vccd1 _28007__473/HI _28007_/A sky130_fd_sc_hd__conb_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17211_ _27082_/Q _27114_/Q _17234_/S vssd1 vssd1 vccd1 vccd1 _17211_/X sky130_fd_sc_hd__mux2_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _15701_/A _14426_/B vssd1 vssd1 vccd1 vccd1 _14423_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26409_ _20737_/X _26409_/D vssd1 vssd1 vccd1 vccd1 _26409_/Q sky130_fd_sc_hd__dfxtp_1
X_18191_ _18188_/X _18190_/X _18216_/S vssd1 vssd1 vccd1 vccd1 _18191_/X sky130_fd_sc_hd__mux2_2
X_27389_ _27392_/CLK _27389_/D vssd1 vssd1 vccd1 vccd1 _27389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17142_ _17291_/A vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__buf_2
XFILLER_129_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14354_ _14354_/A _14363_/B vssd1 vssd1 vccd1 vccd1 _14354_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _27008_/Q _13204_/X _13313_/S vssd1 vssd1 vccd1 vccd1 _13306_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17073_ _25816_/Q _26015_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17073_/X sky130_fd_sc_hd__mux2_1
X_14285_ _14372_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16024_ _16240_/C vssd1 vssd1 vccd1 vccd1 _16252_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13236_ _13236_/A vssd1 vssd1 vccd1 vccd1 _27035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _27046_/Q _13166_/X _13167_/S vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17975_ _17973_/X _17974_/X _18056_/S vssd1 vssd1 vccd1 vccd1 _17975_/X sky130_fd_sc_hd__mux2_1
X_13098_ _27359_/Q _13090_/X _13091_/X _27327_/Q _13097_/X vssd1 vssd1 vccd1 vccd1
+ _14734_/A sky130_fd_sc_hd__a221o_4
XFILLER_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19714_ _19714_/A vssd1 vssd1 vccd1 vccd1 _19714_/X sky130_fd_sc_hd__clkbuf_2
X_16926_ _27484_/Q vssd1 vssd1 vccd1 vccd1 _24206_/A sky130_fd_sc_hd__inv_2
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19645_ _25641_/A vssd1 vssd1 vccd1 vccd1 _25726_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16857_ _16857_/A _16332_/X vssd1 vssd1 vccd1 vccd1 _16858_/A sky130_fd_sc_hd__or2b_1
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _13116_/X _26095_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15809_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19576_ _19640_/A vssd1 vssd1 vccd1 vccd1 _19576_/X sky130_fd_sc_hd__clkbuf_1
X_16788_ _16783_/Y _16611_/B _16776_/A _16787_/X vssd1 vssd1 vccd1 vccd1 _16788_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15739_ _26123_/Q _15734_/X _15727_/X _15738_/Y vssd1 vssd1 vccd1 vccd1 _26123_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18527_ _17897_/X _18522_/X _18524_/X _18526_/X _18489_/X vssd1 vssd1 vccd1 vccd1
+ _18528_/C sky130_fd_sc_hd__a221o_1
XFILLER_34_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18458_ _18458_/A vssd1 vssd1 vccd1 vccd1 _18458_/X sky130_fd_sc_hd__buf_2
XFILLER_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17409_ _27381_/Q vssd1 vssd1 vccd1 vccd1 _24061_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18389_ _18389_/A _18322_/X vssd1 vssd1 vccd1 vccd1 _18389_/X sky130_fd_sc_hd__or2b_1
XFILLER_53_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20420_ _20408_/X _20409_/X _20410_/X _20411_/X _20412_/X _20413_/X vssd1 vssd1 vccd1
+ vccd1 _20421_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20351_ _20351_/A vssd1 vssd1 vccd1 vccd1 _20351_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23070_ _27080_/Q _17721_/X _23070_/S vssd1 vssd1 vccd1 vccd1 _23071_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20282_ _20267_/X _20269_/X _20271_/X _20273_/X _20274_/X _20275_/X vssd1 vssd1 vccd1
+ vccd1 _20283_/A sky130_fd_sc_hd__mux4_1
XFILLER_143_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22021_ _22021_/A vssd1 vssd1 vccd1 vccd1 _22086_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26760_ _21972_/X _26760_/D vssd1 vssd1 vccd1 vccd1 _26760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23972_ _23970_/X _23971_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23972_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25711_ _25705_/X _25706_/X _25707_/X _25708_/X _25709_/X _25710_/X vssd1 vssd1 vccd1
+ vccd1 _25712_/A sky130_fd_sc_hd__mux4_1
X_22923_ _22955_/A vssd1 vssd1 vccd1 vccd1 _22923_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26691_ _21730_/X _26691_/D vssd1 vssd1 vccd1 vccd1 _26691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25642_ _25710_/A vssd1 vssd1 vccd1 vccd1 _25642_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22854_ _22870_/A vssd1 vssd1 vccd1 vccd1 _22854_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21805_ _21793_/X _21794_/X _21795_/X _21796_/X _21797_/X _21798_/X vssd1 vssd1 vccd1
+ vccd1 _21806_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25573_ _25572_/X _25552_/X _25553_/X _24933_/B _25554_/X vssd1 vssd1 vccd1 vccd1
+ _25573_/X sky130_fd_sc_hd__o311a_1
XFILLER_25_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22785_ _22785_/A vssd1 vssd1 vccd1 vccd1 _22785_/X sky130_fd_sc_hd__clkbuf_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27312_ _27312_/CLK _27312_/D vssd1 vssd1 vccd1 vccd1 _27312_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24524_ _24522_/Y _24629_/B _24554_/A vssd1 vssd1 vccd1 vccd1 _24524_/X sky130_fd_sc_hd__o21a_1
X_21736_ _21736_/A vssd1 vssd1 vccd1 vccd1 _21736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27243_ _27261_/CLK _27243_/D vssd1 vssd1 vccd1 vccd1 _27243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24455_ _24455_/A vssd1 vssd1 vccd1 vccd1 _27504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21667_ _21737_/A vssd1 vssd1 vccd1 vccd1 _21667_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23406_ _27759_/Q vssd1 vssd1 vccd1 vccd1 _24750_/A sky130_fd_sc_hd__inv_2
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20618_ _20704_/A vssd1 vssd1 vccd1 vccd1 _20685_/A sky130_fd_sc_hd__clkbuf_2
X_27174_ _27174_/CLK _27174_/D vssd1 vssd1 vccd1 vccd1 _27174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24386_ _24386_/A _24638_/A vssd1 vssd1 vccd1 vccd1 _24387_/A sky130_fd_sc_hd__and2_1
XFILLER_193_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21598_ _21598_/A vssd1 vssd1 vccd1 vccd1 _21598_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26125_ _19755_/X _26125_/D vssd1 vssd1 vccd1 vccd1 _26125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23337_ _27757_/Q _23334_/Y _27244_/Q _24763_/A _23336_/Y vssd1 vssd1 vccd1 vccd1
+ _23337_/X sky130_fd_sc_hd__o221a_1
X_20549_ _20549_/A vssd1 vssd1 vccd1 vccd1 _20549_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14070_ _14335_/A _14070_/B vssd1 vssd1 vccd1 vccd1 _14070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26056_ _26056_/CLK _26056_/D vssd1 vssd1 vccd1 vccd1 _26056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23268_ _27746_/Q vssd1 vssd1 vccd1 vccd1 _23268_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25007_ _25007_/A vssd1 vssd1 vccd1 vccd1 _27675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _13021_/A vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__clkbuf_2
X_22219_ _22213_/X _22214_/X _22215_/X _22216_/X _22217_/X _22218_/X vssd1 vssd1 vccd1
+ vccd1 _22220_/A sky130_fd_sc_hd__mux4_1
XFILLER_133_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23199_ _23199_/A vssd1 vssd1 vccd1 vccd1 _27136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17760_ _27434_/Q vssd1 vssd1 vccd1 vccd1 _17760_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14972_ _15710_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14972_/Y sky130_fd_sc_hd__nor2_1
X_26958_ _22662_/X _26958_/D vssd1 vssd1 vccd1 vccd1 _26958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13923_ _13923_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _13923_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16711_ _16711_/A vssd1 vssd1 vccd1 vccd1 _16711_/Y sky130_fd_sc_hd__inv_2
X_25909_ _25909_/CLK _25909_/D vssd1 vssd1 vccd1 vccd1 _25909_/Q sky130_fd_sc_hd__dfxtp_1
X_17691_ _17691_/A vssd1 vssd1 vccd1 vccd1 _25916_/D sky130_fd_sc_hd__clkbuf_1
X_26889_ _22416_/X _26889_/D vssd1 vssd1 vccd1 vccd1 _26889_/Q sky130_fd_sc_hd__dfxtp_1
X_19430_ _19534_/A _19430_/B vssd1 vssd1 vccd1 vccd1 _19430_/X sky130_fd_sc_hd__or2_1
X_16642_ _16638_/A _16638_/B _16877_/A vssd1 vssd1 vccd1 vccd1 _16642_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _13872_/A vssd1 vssd1 vccd1 vccd1 _13940_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16573_ _16572_/X _16652_/B _16651_/A vssd1 vssd1 vccd1 vccd1 _16573_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19361_ _19350_/X _19355_/X _19359_/X _19290_/X _19360_/X vssd1 vssd1 vccd1 vccd1
+ _19362_/C sky130_fd_sc_hd__a221o_1
X_13785_ _13878_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13785_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18312_ _27812_/Q _26573_/Q _26445_/Q _26125_/Q _18242_/X _18267_/X vssd1 vssd1 vccd1
+ vccd1 _18312_/X sky130_fd_sc_hd__mux4_2
XFILLER_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15524_ _15524_/A vssd1 vssd1 vccd1 vccd1 _26214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19292_ _19362_/A _19292_/B _19292_/C vssd1 vssd1 vccd1 vccd1 _19293_/A sky130_fd_sc_hd__and3_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18243_ _27809_/Q _26570_/Q _26442_/Q _26122_/Q _18242_/X _18126_/X vssd1 vssd1 vccd1
+ vccd1 _18243_/X sky130_fd_sc_hd__mux4_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15455_ _15455_/A vssd1 vssd1 vccd1 vccd1 _26245_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ _14406_/A _14412_/B vssd1 vssd1 vccd1 vccd1 _14406_/Y sky130_fd_sc_hd__nor2_1
XFILLER_198_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18174_ _18172_/X _18173_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18174_/X sky130_fd_sc_hd__mux2_1
X_15386_ _14782_/X _26275_/Q _15390_/S vssd1 vssd1 vccd1 vccd1 _15387_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17125_ _27075_/Q _27107_/Q _17173_/S vssd1 vssd1 vccd1 vccd1 _17125_/X sky130_fd_sc_hd__mux2_1
X_14337_ _14365_/A vssd1 vssd1 vccd1 vccd1 _14337_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17056_ input36/X vssd1 vssd1 vccd1 vccd1 _17181_/A sky130_fd_sc_hd__buf_2
X_14268_ _14356_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14268_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16007_ _16244_/B _16244_/C vssd1 vssd1 vccd1 vccd1 _16136_/A sky130_fd_sc_hd__and2_1
X_13219_ _27274_/Q _13237_/B vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__and2_1
XFILLER_98_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14199_ _14225_/A vssd1 vssd1 vccd1 vccd1 _14199_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater302 _27659_/CLK vssd1 vssd1 vccd1 vccd1 _27649_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17958_ _17779_/X _17953_/X _17957_/X _17932_/X vssd1 vssd1 vccd1 vccd1 _17970_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater313 _27705_/CLK vssd1 vssd1 vccd1 vccd1 _27709_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater324 _27773_/CLK vssd1 vssd1 vccd1 vccd1 _27770_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater335 _27758_/CLK vssd1 vssd1 vccd1 vccd1 _27760_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater346 _27582_/CLK vssd1 vssd1 vccd1 vccd1 _27578_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_111_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16909_ _16908_/A _16908_/B _16087_/X vssd1 vssd1 vccd1 vccd1 _16909_/Y sky130_fd_sc_hd__a21oi_1
Xrepeater357 _27542_/CLK vssd1 vssd1 vccd1 vccd1 _27573_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17889_ _18000_/A vssd1 vssd1 vccd1 vccd1 _18380_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_455 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater368 _27209_/CLK vssd1 vssd1 vccd1 vccd1 _27103_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater379 _27225_/CLK vssd1 vssd1 vccd1 vccd1 _27559_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_81_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19628_ _19628_/A vssd1 vssd1 vccd1 vccd1 _19628_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19559_ _26169_/Q _26105_/Q _27033_/Q _27001_/Q _18930_/A _19482_/X vssd1 vssd1 vccd1
+ vccd1 _19560_/B sky130_fd_sc_hd__mux4_1
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22570_ _22570_/A vssd1 vssd1 vccd1 vccd1 _22570_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21521_ _21513_/X _21514_/X _21515_/X _21516_/X _21517_/X _21518_/X vssd1 vssd1 vccd1
+ vccd1 _21522_/A sky130_fd_sc_hd__mux4_1
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27999__465 vssd1 vssd1 vccd1 vccd1 _27999__465/HI _27999_/A sky130_fd_sc_hd__conb_1
X_24240_ _24240_/A _24250_/B vssd1 vssd1 vccd1 vccd1 _24241_/A sky130_fd_sc_hd__and2_1
X_21452_ _21452_/A vssd1 vssd1 vccd1 vccd1 _21452_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20403_ _20403_/A vssd1 vssd1 vccd1 vccd1 _20403_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21383_ _21373_/X _21374_/X _21375_/X _21376_/X _21377_/X _21378_/X vssd1 vssd1 vccd1
+ vccd1 _21384_/A sky130_fd_sc_hd__mux4_1
X_24171_ _27462_/Q _24173_/B vssd1 vssd1 vccd1 vccd1 _24172_/A sky130_fd_sc_hd__and2_1
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_416 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23122_ _23122_/A vssd1 vssd1 vccd1 vccd1 _27102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20334_ _20334_/A vssd1 vssd1 vccd1 vccd1 _20334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27930_ _27930_/A _15955_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
X_20265_ _20265_/A vssd1 vssd1 vccd1 vccd1 _20265_/X sky130_fd_sc_hd__clkbuf_1
X_23053_ _27072_/Q _17696_/X _23059_/S vssd1 vssd1 vccd1 vccd1 _23054_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22004_ _22072_/A vssd1 vssd1 vccd1 vccd1 _22004_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20196_ _20181_/X _20183_/X _20185_/X _20187_/X _20188_/X _20189_/X vssd1 vssd1 vccd1
+ vccd1 _20197_/A sky130_fd_sc_hd__mux4_1
XFILLER_89_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26812_ _22152_/X _26812_/D vssd1 vssd1 vccd1 vccd1 _26812_/Q sky130_fd_sc_hd__dfxtp_1
X_27792_ _27792_/CLK _27792_/D vssd1 vssd1 vccd1 vccd1 _27982_/A sky130_fd_sc_hd__dfxtp_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26743_ _21908_/X _26743_/D vssd1 vssd1 vccd1 vccd1 _26743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23955_ _24002_/A vssd1 vssd1 vccd1 vccd1 _23955_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22906_ _22906_/A vssd1 vssd1 vccd1 vccd1 _22906_/X sky130_fd_sc_hd__clkbuf_1
X_26674_ _21664_/X _26674_/D vssd1 vssd1 vccd1 vccd1 _26674_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23886_ _23884_/X _23885_/X _23893_/S vssd1 vssd1 vccd1 vccd1 _23886_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25625_ _24987_/S _27982_/A _25625_/S vssd1 vssd1 vccd1 vccd1 _25626_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_447 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22837_ _22869_/A vssd1 vssd1 vccd1 vccd1 _22837_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _26941_/Q _13558_/X _13553_/X _13569_/Y vssd1 vssd1 vccd1 vccd1 _26941_/D
+ sky130_fd_sc_hd__a31o_1
X_25556_ _25530_/X _25274_/B _25555_/X _25543_/X vssd1 vssd1 vccd1 vccd1 _25556_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22768_ _22784_/A vssd1 vssd1 vccd1 vccd1 _22768_/X sky130_fd_sc_hd__clkbuf_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24507_ _27603_/Q _24509_/B vssd1 vssd1 vccd1 vccd1 _24508_/A sky130_fd_sc_hd__and2_1
XFILLER_9_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21719_ _21705_/X _21706_/X _21707_/X _21708_/X _21709_/X _21710_/X vssd1 vssd1 vccd1
+ vccd1 _21720_/A sky130_fd_sc_hd__mux4_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25487_ _25517_/A vssd1 vssd1 vccd1 vccd1 _25487_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22699_ _22699_/A vssd1 vssd1 vccd1 vccd1 _22699_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A vssd1 vssd1 vccd1 vccd1 _26340_/D sky130_fd_sc_hd__clkbuf_1
X_27226_ _27559_/CLK _27226_/D vssd1 vssd1 vccd1 vccd1 _27226_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24438_ _24438_/A vssd1 vssd1 vccd1 vccd1 _27496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27157_ _27157_/CLK _27157_/D vssd1 vssd1 vccd1 vccd1 _27157_/Q sky130_fd_sc_hd__dfxtp_1
X_15171_ _26370_/Q _13395_/X _15173_/S vssd1 vssd1 vccd1 vccd1 _15172_/A sky130_fd_sc_hd__mux2_1
X_24369_ _24369_/A vssd1 vssd1 vccd1 vccd1 _27466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14122_ _26757_/Q _14117_/X _14120_/X _14121_/Y vssd1 vssd1 vccd1 vccd1 _26757_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26108_ _19691_/X _26108_/D vssd1 vssd1 vccd1 vccd1 _26108_/Q sky130_fd_sc_hd__dfxtp_1
X_27088_ _27088_/CLK _27088_/D vssd1 vssd1 vccd1 vccd1 _27088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26039_ _26039_/CLK _26039_/D vssd1 vssd1 vccd1 vccd1 _26039_/Q sky130_fd_sc_hd__dfxtp_1
X_14053_ _14408_/A _14060_/B vssd1 vssd1 vccd1 vccd1 _14053_/Y sky130_fd_sc_hd__nor2_1
X_18930_ _18930_/A vssd1 vssd1 vccd1 vccd1 _18930_/X sky130_fd_sc_hd__buf_4
XFILLER_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _13004_/A vssd1 vssd1 vccd1 vccd1 _27797_/D sky130_fd_sc_hd__clkbuf_1
X_18861_ _18814_/X _18860_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _18861_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17812_ _27595_/Q vssd1 vssd1 vccd1 vccd1 _18156_/A sky130_fd_sc_hd__buf_2
XFILLER_95_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _19297_/A vssd1 vssd1 vccd1 vccd1 _19465_/A sky130_fd_sc_hd__buf_2
X_17743_ _17743_/A vssd1 vssd1 vccd1 vccd1 _25932_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14955_ _14810_/X _26458_/Q _14955_/S vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13906_ _13919_/A vssd1 vssd1 vccd1 vccd1 _13906_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17674_ _24061_/A _17674_/B _17674_/C vssd1 vssd1 vccd1 vccd1 _18691_/A sky130_fd_sc_hd__or3_1
X_14886_ _14942_/A vssd1 vssd1 vccd1 vccd1 _14955_/S sky130_fd_sc_hd__buf_2
XFILLER_36_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19413_ _26962_/Q _26930_/Q _26898_/Q _26866_/Q _19343_/X _19412_/X vssd1 vssd1 vccd1
+ vccd1 _19413_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13837_ _26847_/Q _13832_/X _13833_/X _13836_/Y vssd1 vssd1 vccd1 vccd1 _26847_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16625_ _16625_/A _16625_/B vssd1 vssd1 vccd1 vccd1 _16626_/A sky130_fd_sc_hd__or2_1
XFILLER_189_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19344_ _26959_/Q _26927_/Q _26895_/Q _26863_/Q _19343_/X _19253_/X vssd1 vssd1 vccd1
+ vccd1 _19344_/X sky130_fd_sc_hd__mux4_1
X_16556_ _25969_/Q vssd1 vssd1 vccd1 vccd1 _16556_/Y sky130_fd_sc_hd__inv_2
X_13768_ _13859_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13768_/Y sky130_fd_sc_hd__nor2_1
X_15507_ _15507_/A vssd1 vssd1 vccd1 vccd1 _26222_/D sky130_fd_sc_hd__clkbuf_1
X_19275_ _19273_/X _19274_/X _19229_/X vssd1 vssd1 vccd1 vccd1 _19275_/X sky130_fd_sc_hd__o21a_1
X_16487_ _16809_/A vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13699_ _26898_/Q _13697_/X _13692_/X _13698_/Y vssd1 vssd1 vccd1 vccd1 _26898_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18226_ _17912_/X _18225_/X _17915_/X vssd1 vssd1 vccd1 vccd1 _18226_/X sky130_fd_sc_hd__o21a_1
X_15438_ _26252_/Q _13363_/X _15440_/S vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18157_ _18157_/A _18156_/X vssd1 vssd1 vccd1 vccd1 _18157_/X sky130_fd_sc_hd__or2b_1
XFILLER_157_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15369_/A vssd1 vssd1 vccd1 vccd1 _26283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17108_ _17380_/S vssd1 vssd1 vccd1 vccd1 _17158_/S sky130_fd_sc_hd__clkbuf_2
X_18088_ _17995_/X _18082_/X _18084_/X _18087_/X _18016_/X vssd1 vssd1 vccd1 vccd1
+ _18097_/B sky130_fd_sc_hd__a221o_1
XFILLER_116_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17039_ _17039_/A vssd1 vssd1 vccd1 vccd1 _27918_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20050_ _20044_/X _20045_/X _20046_/X _20047_/X _20048_/X _20049_/X vssd1 vssd1 vccd1
+ vccd1 _20051_/A sky130_fd_sc_hd__mux4_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater110 _27126_/CLK vssd1 vssd1 vccd1 vccd1 _27123_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater121 _27675_/CLK vssd1 vssd1 vccd1 vccd1 _27672_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater132 _27845_/CLK vssd1 vssd1 vccd1 vccd1 _27148_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater143 _27127_/CLK vssd1 vssd1 vccd1 vccd1 _27095_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater154 _27383_/CLK vssd1 vssd1 vccd1 vccd1 _27308_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater165 _27792_/CLK vssd1 vssd1 vccd1 vccd1 _27130_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater176 _27111_/CLK vssd1 vssd1 vccd1 vccd1 _27077_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_27_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23740_ _23849_/A vssd1 vssd1 vccd1 vccd1 _23740_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20952_ _20952_/A vssd1 vssd1 vccd1 vccd1 _20952_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater187 _27415_/CLK vssd1 vssd1 vccd1 vccd1 _27416_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater198 _27826_/CLK vssd1 vssd1 vccd1 vccd1 _26012_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_739 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23671_ _23671_/A vssd1 vssd1 vccd1 vccd1 _27241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _20864_/X _20865_/X _20866_/X _20867_/X _20870_/X _20874_/X vssd1 vssd1 vccd1
+ vccd1 _20884_/A sky130_fd_sc_hd__mux4_1
XFILLER_42_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25410_ _25410_/A vssd1 vssd1 vccd1 vccd1 _27743_/D sky130_fd_sc_hd__clkbuf_1
X_22622_ _22622_/A vssd1 vssd1 vccd1 vccd1 _22622_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26390_ _20675_/X _26390_/D vssd1 vssd1 vccd1 vccd1 _26390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_912 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25341_ _25354_/A _27516_/Q vssd1 vssd1 vccd1 vccd1 _25341_/Y sky130_fd_sc_hd__nand2_1
X_22553_ _22539_/X _22542_/X _22545_/X _22548_/X _22549_/X _22550_/X vssd1 vssd1 vccd1
+ vccd1 _22554_/A sky130_fd_sc_hd__mux4_1
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21504_ _21504_/A vssd1 vssd1 vccd1 vccd1 _21504_/X sky130_fd_sc_hd__clkbuf_1
X_25272_ _25272_/A _25272_/B _25272_/C vssd1 vssd1 vccd1 vccd1 _25273_/B sky130_fd_sc_hd__and3_1
X_22484_ _22484_/A vssd1 vssd1 vccd1 vccd1 _22484_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27011_ _22846_/X _27011_/D vssd1 vssd1 vccd1 vccd1 _27011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24223_ _24298_/A vssd1 vssd1 vccd1 vccd1 _24304_/A sky130_fd_sc_hd__clkbuf_2
X_21435_ _21427_/X _21428_/X _21429_/X _21430_/X _21431_/X _21432_/X vssd1 vssd1 vccd1
+ vccd1 _21436_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24154_ _27454_/Q _24162_/B vssd1 vssd1 vccd1 vccd1 _24155_/A sky130_fd_sc_hd__and2_1
X_21366_ _21366_/A vssd1 vssd1 vccd1 vccd1 _21366_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23105_ _27096_/Q _17772_/X _23107_/S vssd1 vssd1 vccd1 vccd1 _23106_/A sky130_fd_sc_hd__mux2_1
X_20317_ _20317_/A vssd1 vssd1 vccd1 vccd1 _20317_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24085_ _24085_/A vssd1 vssd1 vccd1 vccd1 _27318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21297_ _21285_/X _21286_/X _21287_/X _21288_/X _21289_/X _21290_/X vssd1 vssd1 vccd1
+ vccd1 _21298_/A sky130_fd_sc_hd__mux4_1
XFILLER_116_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23036_ _23109_/A _23182_/B _23109_/C vssd1 vssd1 vccd1 vccd1 _24001_/A sky130_fd_sc_hd__and3_2
XFILLER_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20248_ _20248_/A vssd1 vssd1 vccd1 vccd1 _20248_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27844_ _27844_/CLK _27844_/D vssd1 vssd1 vccd1 vccd1 _27844_/Q sky130_fd_sc_hd__dfxtp_1
X_20179_ _20179_/A vssd1 vssd1 vccd1 vccd1 _20179_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24987_ _24985_/X _24986_/X _24987_/S vssd1 vssd1 vccd1 vccd1 _24987_/X sky130_fd_sc_hd__mux2_1
X_27775_ _27776_/CLK _27775_/D vssd1 vssd1 vccd1 vccd1 _27775_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _14740_/A vssd1 vssd1 vccd1 vccd1 _14740_/X sky130_fd_sc_hd__clkbuf_4
X_26726_ _21856_/X _26726_/D vssd1 vssd1 vccd1 vccd1 _26726_/Q sky130_fd_sc_hd__dfxtp_1
X_23938_ _23936_/X _23937_/X _23938_/S vssd1 vssd1 vccd1 vccd1 _23938_/X sky130_fd_sc_hd__mux2_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26657_ _21610_/X _26657_/D vssd1 vssd1 vccd1 vccd1 _26657_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _14671_/A vssd1 vssd1 vccd1 vccd1 _14671_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23869_ _27077_/Q _27109_/Q _23892_/S vssd1 vssd1 vccd1 vccd1 _23869_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _16774_/A _16410_/B vssd1 vssd1 vccd1 vccd1 _16411_/B sky130_fd_sc_hd__xor2_1
X_13622_ _26925_/Q _13613_/X _13616_/X _13621_/Y vssd1 vssd1 vccd1 vccd1 _26925_/D
+ sky130_fd_sc_hd__a31o_1
X_25608_ _18594_/A _25351_/B _25607_/X _25568_/A vssd1 vssd1 vccd1 vccd1 _25608_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_77_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17390_ _20788_/A vssd1 vssd1 vccd1 vccd1 _25653_/A sky130_fd_sc_hd__buf_6
X_26588_ _21370_/X _26588_/D vssd1 vssd1 vccd1 vccd1 _26588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16341_ _16759_/A _16759_/B vssd1 vssd1 vccd1 vccd1 _16864_/A sky130_fd_sc_hd__or2_1
XFILLER_185_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13553_ _13553_/A vssd1 vssd1 vccd1 vccd1 _13553_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25539_ _25539_/A vssd1 vssd1 vccd1 vccd1 _25539_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater79 _27437_/CLK vssd1 vssd1 vccd1 vccd1 _27430_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19060_ _19060_/A vssd1 vssd1 vccd1 vccd1 _26050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_765 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16272_ _27536_/Q _16254_/S vssd1 vssd1 vccd1 vccd1 _16272_/X sky130_fd_sc_hd__or2b_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13484_ _16289_/A vssd1 vssd1 vccd1 vccd1 _13887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _18011_/A vssd1 vssd1 vccd1 vccd1 _18011_/X sky130_fd_sc_hd__clkbuf_4
X_15223_ _14756_/X _26347_/Q _15223_/S vssd1 vssd1 vccd1 vccd1 _15224_/A sky130_fd_sc_hd__mux2_1
X_27209_ _27209_/CLK _27209_/D vssd1 vssd1 vccd1 vccd1 _27209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1033 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15154_ _26378_/Q _13369_/X _15162_/S vssd1 vssd1 vccd1 vccd1 _15155_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14105_ _14369_/A _14112_/B vssd1 vssd1 vccd1 vccd1 _14105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15085_ _15085_/A vssd1 vssd1 vccd1 vccd1 _26409_/D sky130_fd_sc_hd__clkbuf_1
X_19962_ _19956_/X _19957_/X _19958_/X _19959_/X _19960_/X _19961_/X vssd1 vssd1 vccd1
+ vccd1 _19963_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14036_ _14396_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14036_/Y sky130_fd_sc_hd__nor2_1
X_18913_ _18913_/A vssd1 vssd1 vccd1 vccd1 _18913_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19893_ _19893_/A vssd1 vssd1 vccd1 vccd1 _19893_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18844_ _18844_/A vssd1 vssd1 vccd1 vccd1 _18989_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18775_ _19553_/S vssd1 vssd1 vccd1 vccd1 _18775_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15987_ _15988_/A vssd1 vssd1 vccd1 vccd1 _15987_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17726_ _25927_/Q _17724_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17727_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14938_ _14785_/X _26466_/Q _14940_/S vssd1 vssd1 vccd1 vccd1 _14939_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17657_ _17657_/A vssd1 vssd1 vccd1 vccd1 _25899_/D sky130_fd_sc_hd__clkbuf_1
X_14869_ _14869_/A vssd1 vssd1 vccd1 vccd1 _26497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _16692_/A _16692_/B _16692_/C vssd1 vssd1 vccd1 vccd1 _16609_/B sky130_fd_sc_hd__o21ai_1
X_17588_ _17588_/A vssd1 vssd1 vccd1 vccd1 _25868_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19327_ _26158_/Q _26094_/Q _27022_/Q _26990_/Q _19326_/X _19188_/X vssd1 vssd1 vccd1
+ vccd1 _19328_/B sky130_fd_sc_hd__mux4_1
XFILLER_188_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16539_ _16292_/B _16292_/C _16486_/A vssd1 vssd1 vccd1 vccd1 _16540_/B sky130_fd_sc_hd__o21a_1
XFILLER_188_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19258_ _19393_/A vssd1 vssd1 vccd1 vccd1 _19258_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18209_ _18324_/A vssd1 vssd1 vccd1 vccd1 _18209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19189_ _26152_/Q _26088_/Q _27016_/Q _26984_/Q _19165_/X _19188_/X vssd1 vssd1 vccd1
+ vccd1 _19190_/B sky130_fd_sc_hd__mux4_1
XFILLER_145_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21220_ _21220_/A vssd1 vssd1 vccd1 vccd1 _21220_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21151_ _21199_/A vssd1 vssd1 vccd1 vccd1 _21151_/X sky130_fd_sc_hd__clkbuf_2
X_20102_ _20150_/A vssd1 vssd1 vccd1 vccd1 _20102_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21082_ _21114_/A vssd1 vssd1 vccd1 vccd1 _21082_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24910_ _27772_/Q _27771_/Q _24910_/C vssd1 vssd1 vccd1 vccd1 _24918_/B sky130_fd_sc_hd__and3_1
X_20033_ _20065_/A vssd1 vssd1 vccd1 vccd1 _20033_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_923 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25890_ _27145_/CLK _25890_/D vssd1 vssd1 vccd1 vccd1 _25890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24841_ _24841_/A vssd1 vssd1 vccd1 vccd1 _24935_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27560_ _27562_/CLK _27560_/D vssd1 vssd1 vccd1 vccd1 _27560_/Q sky130_fd_sc_hd__dfxtp_1
X_24772_ _24772_/A _24772_/B vssd1 vssd1 vccd1 vccd1 _24772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21984_ _22000_/A vssd1 vssd1 vccd1 vccd1 _21984_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26511_ _21102_/X _26511_/D vssd1 vssd1 vccd1 vccd1 _26511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23723_ _24186_/A vssd1 vssd1 vccd1 vccd1 _24063_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20935_ _20921_/X _20922_/X _20923_/X _20924_/X _20925_/X _20926_/X vssd1 vssd1 vccd1
+ vccd1 _20936_/A sky130_fd_sc_hd__mux4_1
X_27491_ _27534_/CLK _27491_/D vssd1 vssd1 vccd1 vccd1 _27491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26442_ _20859_/X _26442_/D vssd1 vssd1 vccd1 vccd1 _26442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23654_ _23654_/A vssd1 vssd1 vccd1 vccd1 _27233_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _20866_/A vssd1 vssd1 vccd1 vccd1 _20866_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22605_ _22593_/X _22594_/X _22595_/X _22596_/X _22597_/X _22598_/X vssd1 vssd1 vccd1
+ vccd1 _22606_/A sky130_fd_sc_hd__mux4_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26373_ _20613_/X _26373_/D vssd1 vssd1 vccd1 vccd1 _26373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23585_ _24925_/B _27216_/Q _23595_/S vssd1 vssd1 vccd1 vccd1 _23586_/B sky130_fd_sc_hd__mux2_1
X_20797_ _22543_/A vssd1 vssd1 vccd1 vccd1 _21147_/A sky130_fd_sc_hd__clkbuf_2
X_25324_ _25354_/A _27513_/Q _25320_/A vssd1 vssd1 vccd1 vccd1 _25325_/B sky130_fd_sc_hd__a21o_1
XFILLER_167_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22536_ _22536_/A vssd1 vssd1 vccd1 vccd1 _22536_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25255_ _27707_/Q _25223_/X _25253_/Y _25254_/X vssd1 vssd1 vccd1 vccd1 _27707_/D
+ sky130_fd_sc_hd__o211a_1
X_22467_ _22452_/X _22454_/X _22456_/X _22458_/X _22459_/X _22460_/X vssd1 vssd1 vccd1
+ vccd1 _22468_/A sky130_fd_sc_hd__mux4_1
XFILLER_136_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24206_ _24206_/A _24210_/B vssd1 vssd1 vccd1 vccd1 _27370_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21418_ _21418_/A vssd1 vssd1 vccd1 vccd1 _21418_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25186_ _27529_/Q _27497_/Q vssd1 vssd1 vccd1 vccd1 _25188_/A sky130_fd_sc_hd__and2_1
X_22398_ _22398_/A vssd1 vssd1 vccd1 vccd1 _22398_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_185_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24137_ _24137_/A vssd1 vssd1 vccd1 vccd1 _27341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21349_ _21341_/X _21342_/X _21343_/X _21344_/X _21345_/X _21346_/X vssd1 vssd1 vccd1
+ vccd1 _21350_/A sky130_fd_sc_hd__mux4_1
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24068_ _27384_/Q _24072_/B vssd1 vssd1 vccd1 vccd1 _24069_/A sky130_fd_sc_hd__and2_1
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15910_ _15912_/A vssd1 vssd1 vccd1 vccd1 _15910_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23019_ _23009_/X _23010_/X _23011_/X _23012_/X _23013_/X _23014_/X vssd1 vssd1 vccd1
+ vccd1 _23020_/A sky130_fd_sc_hd__mux4_1
XFILLER_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16890_ _16890_/A _16890_/B _16890_/C vssd1 vssd1 vccd1 vccd1 _16890_/X sky130_fd_sc_hd__and3_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _13204_/X _26080_/Q _15849_/S vssd1 vssd1 vccd1 vccd1 _15842_/A sky130_fd_sc_hd__mux2_1
X_27827_ _27827_/CLK _27827_/D vssd1 vssd1 vccd1 vccd1 _27827_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18560_ _26552_/Q _26520_/Q _26488_/Q _27064_/Q _17846_/X _17848_/X vssd1 vssd1 vccd1
+ vccd1 _18560_/X sky130_fd_sc_hd__mux4_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _26110_/Q _15760_/X _15766_/X _15771_/Y vssd1 vssd1 vccd1 vccd1 _26110_/D
+ sky130_fd_sc_hd__a31o_1
X_12984_ _12984_/A vssd1 vssd1 vccd1 vccd1 _27806_/D sky130_fd_sc_hd__clkbuf_1
X_27758_ _27758_/CLK _27758_/D vssd1 vssd1 vccd1 vccd1 _27758_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17511_ _27435_/Q vssd1 vssd1 vccd1 vccd1 _17511_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26709_ _21792_/X _26709_/D vssd1 vssd1 vccd1 vccd1 _26709_/Q sky130_fd_sc_hd__dfxtp_1
X_14723_ _14723_/A vssd1 vssd1 vccd1 vccd1 _26550_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _18509_/A _18491_/B _18491_/C vssd1 vssd1 vccd1 vccd1 _18492_/A sky130_fd_sc_hd__and3_1
XFILLER_18_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27689_ _27693_/CLK _27689_/D vssd1 vssd1 vccd1 vccd1 _27689_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14654_ _15728_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14654_/Y sky130_fd_sc_hd__nor2_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _17440_/X _25816_/Q _17454_/S vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__mux2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _26932_/Q _13599_/X _13603_/X _13604_/Y vssd1 vssd1 vccd1 vccd1 _26932_/D
+ sky130_fd_sc_hd__a31o_1
X_14585_ _26600_/Q _14576_/X _14579_/X _14584_/Y vssd1 vssd1 vccd1 vccd1 _26600_/D
+ sky130_fd_sc_hd__a31o_1
X_17373_ _16992_/X _17372_/X _17342_/X vssd1 vssd1 vccd1 vccd1 _17373_/X sky130_fd_sc_hd__a21bo_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19112_ _26821_/Q _26789_/Q _26757_/Q _26725_/Q _19039_/X _19111_/X vssd1 vssd1 vccd1
+ vccd1 _19113_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16324_ _14801_/A _16501_/A _16412_/A _25947_/Q _16323_/Y vssd1 vssd1 vccd1 vccd1
+ _16752_/B sky130_fd_sc_hd__a221o_1
X_13536_ _27345_/Q _13529_/X _13530_/X _27313_/Q _13176_/X vssd1 vssd1 vccd1 vccd1
+ _14497_/A sky130_fd_sc_hd__a221oi_4
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19043_ _18996_/X _19042_/X _18941_/X vssd1 vssd1 vccd1 vccd1 _19043_/X sky130_fd_sc_hd__o21a_1
X_16255_ _16459_/A _16453_/A vssd1 vssd1 vccd1 vccd1 _16255_/Y sky130_fd_sc_hd__nor2_1
XFILLER_199_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ _13876_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13467_/Y sky130_fd_sc_hd__nor2_1
XFILLER_199_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _14731_/X _26355_/Q _15212_/S vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16186_ _27519_/Q _27576_/Q vssd1 vssd1 vccd1 vccd1 _16186_/X sky130_fd_sc_hd__or2b_1
X_13398_ _16206_/A vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__clkbuf_4
X_15137_ _15137_/A vssd1 vssd1 vccd1 vccd1 _26386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19945_ _19977_/A vssd1 vssd1 vccd1 vccd1 _19945_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15068_ _14740_/X _26416_/Q _15068_/S vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14019_ _14038_/A vssd1 vssd1 vccd1 vccd1 _14019_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19876_ _19866_/X _19867_/X _19868_/X _19869_/X _19870_/X _19871_/X vssd1 vssd1 vccd1
+ vccd1 _19877_/A sky130_fd_sc_hd__mux4_1
X_18827_ _26394_/Q _26362_/Q _26330_/Q _26298_/Q _18824_/X _18826_/X vssd1 vssd1 vccd1
+ vccd1 _18827_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18758_ _18758_/A vssd1 vssd1 vccd1 vccd1 _26039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17709_ _17776_/S vssd1 vssd1 vccd1 vccd1 _17722_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18689_ _26009_/Q _17775_/X _18689_/S vssd1 vssd1 vccd1 vccd1 _18690_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20720_ _20703_/X _20705_/X _20707_/X _20709_/X _20710_/X _20711_/X vssd1 vssd1 vccd1
+ vccd1 _20721_/A sky130_fd_sc_hd__mux4_1
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20651_ _20651_/A vssd1 vssd1 vccd1 vccd1 _20651_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23370_ _27770_/Q vssd1 vssd1 vccd1 vccd1 _24778_/A sky130_fd_sc_hd__inv_2
X_20582_ _20598_/A vssd1 vssd1 vccd1 vccd1 _20582_/X sky130_fd_sc_hd__clkbuf_1
X_22321_ _22315_/X _22316_/X _22317_/X _22318_/X _22319_/X _22320_/X vssd1 vssd1 vccd1
+ vccd1 _22322_/A sky130_fd_sc_hd__mux4_1
XFILLER_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25040_ _27232_/Q vssd1 vssd1 vccd1 vccd1 _25074_/S sky130_fd_sc_hd__buf_2
X_22252_ _22252_/A vssd1 vssd1 vccd1 vccd1 _22252_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21203_ _21195_/X _21196_/X _21197_/X _21198_/X _21199_/X _21200_/X vssd1 vssd1 vccd1
+ vccd1 _21204_/A sky130_fd_sc_hd__mux4_1
X_22183_ _22173_/X _22174_/X _22175_/X _22176_/X _22179_/X _22182_/X vssd1 vssd1 vccd1
+ vccd1 _22184_/A sky130_fd_sc_hd__mux4_1
XFILLER_160_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21134_ _21134_/A vssd1 vssd1 vccd1 vccd1 _21134_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26991_ _22776_/X _26991_/D vssd1 vssd1 vccd1 vccd1 _26991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25942_ _27857_/CLK _25942_/D vssd1 vssd1 vccd1 vccd1 _25942_/Q sky130_fd_sc_hd__dfxtp_1
X_21065_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21065_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20016_ _20064_/A vssd1 vssd1 vccd1 vccd1 _20016_/X sky130_fd_sc_hd__clkbuf_2
X_25873_ _27160_/CLK _25873_/D vssd1 vssd1 vccd1 vccd1 _25873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27612_ _27612_/CLK _27612_/D vssd1 vssd1 vccd1 vccd1 _27612_/Q sky130_fd_sc_hd__dfxtp_1
X_24824_ _27640_/Q _24813_/X _24823_/Y _24817_/X vssd1 vssd1 vccd1 vccd1 _27640_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24755_ _27616_/Q _24742_/X _24754_/Y _24746_/X vssd1 vssd1 vccd1 vccd1 _27616_/D
+ sky130_fd_sc_hd__o211a_1
X_27543_ _27582_/CLK _27543_/D vssd1 vssd1 vccd1 vccd1 _27543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ _21999_/A vssd1 vssd1 vccd1 vccd1 _21967_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23706_ _23706_/A vssd1 vssd1 vccd1 vccd1 _27257_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27474_ _27475_/CLK _27474_/D vssd1 vssd1 vccd1 vccd1 _27474_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20918_ _20918_/A vssd1 vssd1 vccd1 vccd1 _20918_/X sky130_fd_sc_hd__clkbuf_1
X_24686_ _16979_/A _24673_/X _24685_/X _24677_/X vssd1 vssd1 vccd1 vccd1 _27592_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21898_ _21914_/A vssd1 vssd1 vccd1 vccd1 _21898_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23637_ _25035_/A vssd1 vssd1 vccd1 vccd1 _23638_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_26425_ _20807_/X _26425_/D vssd1 vssd1 vccd1 vccd1 _26425_/Q sky130_fd_sc_hd__dfxtp_1
X_20849_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20849_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14370_ _26667_/Q _14365_/X _14358_/X _14369_/Y vssd1 vssd1 vccd1 vccd1 _26667_/D
+ sky130_fd_sc_hd__a31o_1
X_26356_ _20559_/X _26356_/D vssd1 vssd1 vccd1 vccd1 _26356_/Q sky130_fd_sc_hd__dfxtp_1
X_23568_ _23577_/A _23568_/B vssd1 vssd1 vccd1 vccd1 _23569_/A sky130_fd_sc_hd__and2_1
XFILLER_70_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25307_ _27713_/Q _25263_/X _25306_/Y _25297_/X vssd1 vssd1 vccd1 vccd1 _27713_/D
+ sky130_fd_sc_hd__o211a_1
X_13321_ _13402_/A vssd1 vssd1 vccd1 vccd1 _13421_/S sky130_fd_sc_hd__buf_2
X_22519_ _22519_/A vssd1 vssd1 vccd1 vccd1 _22519_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26287_ _20313_/X _26287_/D vssd1 vssd1 vccd1 vccd1 _26287_/Q sky130_fd_sc_hd__dfxtp_1
X_23499_ input32/X _23429_/A _23497_/X _23498_/X vssd1 vssd1 vccd1 vccd1 _27192_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _27475_/Q _27371_/Q vssd1 vssd1 vccd1 vccd1 _16040_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_183_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25238_ _27705_/Q _25223_/X _25237_/Y _25214_/X vssd1 vssd1 vccd1 vccd1 _27705_/D
+ sky130_fd_sc_hd__o211a_1
X_13252_ _27032_/Q _13058_/X _13258_/S vssd1 vssd1 vccd1 vccd1 _13253_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25169_ _27527_/Q _27495_/Q vssd1 vssd1 vccd1 vccd1 _25169_/Y sky130_fd_sc_hd__nand2_1
X_13183_ _27344_/Q _13017_/A _13025_/A _27312_/Q _13182_/X vssd1 vssd1 vccd1 vccd1
+ _16235_/A sky130_fd_sc_hd__a221o_4
XFILLER_123_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_630 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17991_ _17983_/X _17985_/X _17989_/X _17854_/X _17990_/X vssd1 vssd1 vccd1 vccd1
+ _17992_/C sky130_fd_sc_hd__a221o_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19730_ _25725_/A vssd1 vssd1 vccd1 vccd1 _19800_/A sky130_fd_sc_hd__clkbuf_2
X_16942_ _27599_/Q _24207_/A _24209_/A _27601_/Q vssd1 vssd1 vccd1 vccd1 _16942_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19661_ _19727_/A vssd1 vssd1 vccd1 vccd1 _19661_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16873_ _24233_/A _24228_/A _24225_/A _16873_/D vssd1 vssd1 vccd1 vccd1 _16874_/D
+ sky130_fd_sc_hd__and4bb_1
X_18612_ _18610_/X _18612_/B vssd1 vssd1 vccd1 vccd1 _18613_/B sky130_fd_sc_hd__and2b_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15824_ _15824_/A vssd1 vssd1 vccd1 vccd1 _26088_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ _19640_/A vssd1 vssd1 vccd1 vccd1 _19592_/X sky130_fd_sc_hd__clkbuf_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18543_ _26423_/Q _26391_/Q _26359_/Q _26327_/Q _18462_/X _18486_/X vssd1 vssd1 vccd1
+ vccd1 _18543_/X sky130_fd_sc_hd__mux4_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ _26117_/Q _15747_/X _15753_/X _15754_/Y vssd1 vssd1 vccd1 vccd1 _26117_/D
+ sky130_fd_sc_hd__a31o_1
X_12967_ _13000_/A vssd1 vssd1 vccd1 vccd1 _12976_/B sky130_fd_sc_hd__clkbuf_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _26555_/Q _14698_/X _14631_/B _14705_/Y vssd1 vssd1 vccd1 vccd1 _26555_/D
+ sky130_fd_sc_hd__a31o_1
X_18474_ _18474_/A vssd1 vssd1 vccd1 vccd1 _18474_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_360 _25583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15686_ _15686_/A vssd1 vssd1 vccd1 vccd1 _26142_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17425_ _17524_/S vssd1 vssd1 vccd1 vccd1 _17438_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_382 _13389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14637_ _15710_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ _17354_/X _17355_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17356_/X sky130_fd_sc_hd__mux2_2
X_14568_ _26607_/Q _14563_/X _14566_/X _14567_/Y vssd1 vssd1 vccd1 vccd1 _26607_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16307_ _16308_/A _16308_/B vssd1 vssd1 vccd1 vccd1 _16309_/A sky130_fd_sc_hd__nand2_1
X_13519_ _27348_/Q _13019_/A _13027_/A _27316_/Q _13159_/X vssd1 vssd1 vccd1 vccd1
+ _16243_/A sky130_fd_sc_hd__a221oi_4
XFILLER_173_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14499_ _26628_/Q _14496_/X _14492_/X _14498_/Y vssd1 vssd1 vccd1 vccd1 _26628_/D
+ sky130_fd_sc_hd__a31o_1
X_17287_ _17287_/A vssd1 vssd1 vccd1 vccd1 _27938_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19026_ _26145_/Q _26081_/Q _27009_/Q _26977_/Q _18882_/X _18950_/X vssd1 vssd1 vccd1
+ vccd1 _19027_/B sky130_fd_sc_hd__mux4_1
X_16238_ _16408_/A _16406_/A vssd1 vssd1 vccd1 vccd1 _16447_/D sky130_fd_sc_hd__or2_1
XFILLER_162_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16169_ _16169_/A _16249_/B _16240_/C vssd1 vssd1 vccd1 vccd1 _16169_/X sky130_fd_sc_hd__and3_1
XFILLER_173_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19928_ _19976_/A vssd1 vssd1 vccd1 vccd1 _19928_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19859_ _19859_/A vssd1 vssd1 vccd1 vccd1 _19859_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22870_ _22870_/A vssd1 vssd1 vccd1 vccd1 _22870_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21821_ _21809_/X _21810_/X _21811_/X _21812_/X _21813_/X _21814_/X vssd1 vssd1 vccd1
+ vccd1 _21822_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24540_ _24552_/A _24540_/B vssd1 vssd1 vccd1 vccd1 _24541_/A sky130_fd_sc_hd__and2_1
X_21752_ _21752_/A vssd1 vssd1 vccd1 vccd1 _21752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20703_ _20770_/A vssd1 vssd1 vccd1 vccd1 _20703_/X sky130_fd_sc_hd__clkbuf_1
X_24471_ _24471_/A vssd1 vssd1 vccd1 vccd1 _27511_/D sky130_fd_sc_hd__clkbuf_1
X_21683_ _21667_/X _21670_/X _21673_/X _21676_/X _21677_/X _21678_/X vssd1 vssd1 vccd1
+ vccd1 _21684_/A sky130_fd_sc_hd__mux4_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26210_ _20051_/X _26210_/D vssd1 vssd1 vccd1 vccd1 _26210_/Q sky130_fd_sc_hd__dfxtp_1
X_23422_ input9/X _23415_/X _23419_/X _23421_/X vssd1 vssd1 vccd1 vccd1 _27162_/D
+ sky130_fd_sc_hd__o211a_1
X_27190_ _27190_/CLK _27190_/D vssd1 vssd1 vccd1 vccd1 _27190_/Q sky130_fd_sc_hd__dfxtp_1
X_20634_ _20617_/X _20619_/X _20621_/X _20623_/X _20624_/X _20625_/X vssd1 vssd1 vccd1
+ vccd1 _20635_/A sky130_fd_sc_hd__mux4_1
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26141_ _19805_/X _26141_/D vssd1 vssd1 vccd1 vccd1 _26141_/Q sky130_fd_sc_hd__dfxtp_1
X_23353_ _27775_/Q vssd1 vssd1 vccd1 vccd1 _24925_/A sky130_fd_sc_hd__buf_4
X_20565_ _20565_/A vssd1 vssd1 vccd1 vccd1 _20565_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22304_ _22336_/A vssd1 vssd1 vccd1 vccd1 _22304_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26072_ _27332_/CLK _26072_/D vssd1 vssd1 vccd1 vccd1 _26072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23284_ input43/X vssd1 vssd1 vccd1 vccd1 _23284_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20496_ _20512_/A vssd1 vssd1 vccd1 vccd1 _20496_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_672 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25023_ _25021_/X _25022_/X _25031_/S vssd1 vssd1 vccd1 vccd1 _25023_/X sky130_fd_sc_hd__mux2_1
X_22235_ _22229_/X _22230_/X _22231_/X _22232_/X _22233_/X _22234_/X vssd1 vssd1 vccd1
+ vccd1 _22236_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22166_ _22166_/A vssd1 vssd1 vccd1 vccd1 _22166_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21117_ _21109_/X _21110_/X _21111_/X _21112_/X _21113_/X _21114_/X vssd1 vssd1 vccd1
+ vccd1 _21118_/A sky130_fd_sc_hd__mux4_1
XFILLER_121_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22097_ _22083_/X _22084_/X _22085_/X _22086_/X _22088_/X _22090_/X vssd1 vssd1 vccd1
+ vccd1 _22098_/A sky130_fd_sc_hd__mux4_1
X_26974_ _22714_/X _26974_/D vssd1 vssd1 vccd1 vccd1 _26974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25925_ _25925_/CLK _25925_/D vssd1 vssd1 vccd1 vccd1 _25925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21048_ _21048_/A vssd1 vssd1 vccd1 vccd1 _21048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _13870_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25856_ _25925_/CLK _25856_/D vssd1 vssd1 vccd1 vccd1 _25856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24807_ _27635_/Q _24798_/X _24806_/Y _24801_/X vssd1 vssd1 vccd1 vccd1 _27635_/D
+ sky130_fd_sc_hd__o211a_1
X_25787_ _25787_/A vssd1 vssd1 vccd1 vccd1 _27848_/D sky130_fd_sc_hd__clkbuf_1
X_22999_ _22993_/X _22994_/X _22995_/X _22996_/X _22997_/X _22998_/X vssd1 vssd1 vccd1
+ vccd1 _23000_/A sky130_fd_sc_hd__mux4_1
X_27526_ _27527_/CLK _27526_/D vssd1 vssd1 vccd1 vccd1 _27526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _15540_/A vssd1 vssd1 vccd1 vccd1 _26207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24738_ _27611_/Q _24727_/X _24737_/Y _24729_/X vssd1 vssd1 vccd1 vccd1 _27611_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _26237_/Q _13411_/X _15473_/S vssd1 vssd1 vccd1 vccd1 _15472_/A sky130_fd_sc_hd__mux2_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27457_ _27458_/CLK _27457_/D vssd1 vssd1 vccd1 vccd1 _27457_/Q sky130_fd_sc_hd__dfxtp_1
X_24669_ _27170_/Q _24671_/B vssd1 vssd1 vccd1 vccd1 _24669_/X sky130_fd_sc_hd__or2_1
XFILLER_188_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17177_/X _17204_/X _17207_/X _17209_/X vssd1 vssd1 vccd1 vccd1 _17210_/X
+ sky130_fd_sc_hd__o22a_1
X_14422_ _16099_/A vssd1 vssd1 vccd1 vccd1 _15701_/A sky130_fd_sc_hd__buf_2
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26408_ _20735_/X _26408_/D vssd1 vssd1 vccd1 vccd1 _26408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18190_ _26407_/Q _26375_/Q _26343_/Q _26311_/Q _18189_/X _18073_/X vssd1 vssd1 vccd1
+ vccd1 _18190_/X sky130_fd_sc_hd__mux4_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27388_ _27388_/CLK _27388_/D vssd1 vssd1 vccd1 vccd1 _27388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14353_ _14393_/A vssd1 vssd1 vccd1 vccd1 _14363_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17141_ _17141_/A vssd1 vssd1 vccd1 vccd1 _27926_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_156_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26339_ _20495_/X _26339_/D vssd1 vssd1 vccd1 vccd1 _26339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13304_ _13304_/A vssd1 vssd1 vccd1 vccd1 _13313_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_156_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17072_ _17029_/X _17072_/B vssd1 vssd1 vccd1 vccd1 _17072_/X sky130_fd_sc_hd__and2b_1
X_14284_ _14311_/A vssd1 vssd1 vccd1 vccd1 _14284_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13235_ _27035_/Q _13234_/X _13241_/S vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__mux2_1
X_16023_ _16197_/C vssd1 vssd1 vccd1 vccd1 _16240_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_28009_ _28009_/A _15918_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
XFILLER_156_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ _16240_/A vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17974_ _26943_/Q _26911_/Q _26879_/Q _26847_/Q _17922_/X _17951_/X vssd1 vssd1 vccd1
+ vccd1 _17974_/X sky130_fd_sc_hd__mux4_2
X_13097_ _27295_/Q _13109_/B vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__and2_2
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19713_ _19729_/A vssd1 vssd1 vccd1 vccd1 _19713_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16925_ _27485_/Q vssd1 vssd1 vccd1 vccd1 _24207_/A sky130_fd_sc_hd__inv_2
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19644_ _19714_/A vssd1 vssd1 vccd1 vccd1 _19644_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16856_ _16852_/Y _16853_/X _16855_/X vssd1 vssd1 vccd1 vccd1 _25617_/A sky130_fd_sc_hd__a21oi_2
XFILLER_168_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _15853_/S vssd1 vssd1 vccd1 vccd1 _15816_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19575_ _19836_/A vssd1 vssd1 vccd1 vccd1 _19640_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16787_ _16446_/Y _16479_/A _16785_/Y _16786_/X vssd1 vssd1 vccd1 vccd1 _16787_/X
+ sky130_fd_sc_hd__o211a_1
X_13999_ _14369_/A _14010_/B vssd1 vssd1 vccd1 vccd1 _13999_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18526_ _17827_/X _18525_/X _17838_/X vssd1 vssd1 vccd1 vccd1 _18526_/X sky130_fd_sc_hd__o21a_1
X_15738_ _15738_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15738_/Y sky130_fd_sc_hd__nor2_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _18457_/A _18322_/X vssd1 vssd1 vccd1 vccd1 _18457_/X sky130_fd_sc_hd__or2b_1
XFILLER_179_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15669_ _15680_/A vssd1 vssd1 vccd1 vccd1 _15678_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_190 _16451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17408_ _27408_/Q vssd1 vssd1 vccd1 vccd1 _17408_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18388_ _26160_/Q _26096_/Q _27024_/Q _26992_/Q _18298_/X _18387_/X vssd1 vssd1 vccd1
+ vccd1 _18389_/A sky130_fd_sc_hd__mux4_1
XFILLER_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17339_ _25939_/Q _26005_/Q _17370_/S vssd1 vssd1 vccd1 vccd1 _17340_/B sky130_fd_sc_hd__mux2_1
XFILLER_179_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20350_ _20334_/X _20335_/X _20336_/X _20337_/X _20339_/X _20341_/X vssd1 vssd1 vccd1
+ vccd1 _20351_/A sky130_fd_sc_hd__mux4_1
XFILLER_101_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19009_ _19007_/X _19008_/X _19057_/S vssd1 vssd1 vccd1 vccd1 _19009_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20281_ _20281_/A vssd1 vssd1 vccd1 vccd1 _20281_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22020_ _22085_/A vssd1 vssd1 vccd1 vccd1 _22020_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23971_ _27088_/Q _27120_/Q _23986_/S vssd1 vssd1 vccd1 vccd1 _23971_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22922_ _22922_/A vssd1 vssd1 vccd1 vccd1 _22922_/X sky130_fd_sc_hd__clkbuf_1
X_25710_ _25710_/A vssd1 vssd1 vccd1 vccd1 _25710_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26690_ _21728_/X _26690_/D vssd1 vssd1 vccd1 vccd1 _26690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22853_ _22869_/A vssd1 vssd1 vccd1 vccd1 _22853_/X sky130_fd_sc_hd__clkbuf_1
X_25641_ _25641_/A vssd1 vssd1 vccd1 vccd1 _25710_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21804_ _21804_/A vssd1 vssd1 vccd1 vccd1 _21804_/X sky130_fd_sc_hd__clkbuf_1
X_25572_ _25572_/A vssd1 vssd1 vccd1 vccd1 _25572_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22784_ _22784_/A vssd1 vssd1 vccd1 vccd1 _22784_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24523_ _27609_/Q vssd1 vssd1 vccd1 vccd1 _24554_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_27311_ _27311_/CLK _27311_/D vssd1 vssd1 vccd1 vccd1 _27311_/Q sky130_fd_sc_hd__dfxtp_1
X_21735_ _21721_/X _21722_/X _21723_/X _21724_/X _21725_/X _21726_/X vssd1 vssd1 vccd1
+ vccd1 _21736_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24454_ _27625_/Q _24456_/B vssd1 vssd1 vccd1 vccd1 _24455_/A sky130_fd_sc_hd__and2_1
X_27242_ _27258_/CLK _27242_/D vssd1 vssd1 vccd1 vccd1 _27242_/Q sky130_fd_sc_hd__dfxtp_1
X_21666_ _22015_/A vssd1 vssd1 vccd1 vccd1 _21737_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23405_ _27239_/Q vssd1 vssd1 vccd1 vccd1 _23405_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20617_ _20684_/A vssd1 vssd1 vccd1 vccd1 _20617_/X sky130_fd_sc_hd__clkbuf_1
X_27173_ _27593_/CLK _27173_/D vssd1 vssd1 vccd1 vccd1 _27173_/Q sky130_fd_sc_hd__dfxtp_1
X_24385_ _24435_/A vssd1 vssd1 vccd1 vccd1 _24638_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21597_ _21580_/X _21582_/X _21584_/X _21586_/X _21587_/X _21588_/X vssd1 vssd1 vccd1
+ vccd1 _21598_/A sky130_fd_sc_hd__mux4_1
X_26124_ _19743_/X _26124_/D vssd1 vssd1 vccd1 vccd1 _26124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23336_ _27783_/Q _27263_/Q vssd1 vssd1 vccd1 vccd1 _23336_/Y sky130_fd_sc_hd__xnor2_1
X_20548_ _20531_/X _20533_/X _20535_/X _20537_/X _20538_/X _20539_/X vssd1 vssd1 vccd1
+ vccd1 _20549_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26055_ _27325_/CLK _26055_/D vssd1 vssd1 vccd1 vccd1 _26055_/Q sky130_fd_sc_hd__dfxtp_1
X_23267_ input45/X vssd1 vssd1 vccd1 vccd1 _23267_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20479_ _20479_/A vssd1 vssd1 vccd1 vccd1 _20479_/X sky130_fd_sc_hd__clkbuf_1
X_25006_ _27966_/A _25005_/X _25024_/S vssd1 vssd1 vccd1 vccd1 _25007_/A sky130_fd_sc_hd__mux2_1
X_13020_ _13108_/A vssd1 vssd1 vccd1 vccd1 _13021_/A sky130_fd_sc_hd__clkbuf_4
X_22218_ _22250_/A vssd1 vssd1 vccd1 vccd1 _22218_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23198_ _17444_/X _27136_/Q _23204_/S vssd1 vssd1 vccd1 vccd1 _23199_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22149_ _22141_/X _22142_/X _22143_/X _22144_/X _22145_/X _22146_/X vssd1 vssd1 vccd1
+ vccd1 _22150_/A sky130_fd_sc_hd__mux4_1
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26957_ _22660_/X _26957_/D vssd1 vssd1 vccd1 vccd1 _26957_/Q sky130_fd_sc_hd__dfxtp_1
X_14971_ _26454_/Q _14957_/X _14960_/X _14970_/Y vssd1 vssd1 vccd1 vccd1 _26454_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16710_ _16710_/A _16710_/B vssd1 vssd1 vccd1 vccd1 _16710_/X sky130_fd_sc_hd__xor2_1
X_13922_ _26818_/Q _13919_/X _13912_/X _13921_/Y vssd1 vssd1 vccd1 vccd1 _26818_/D
+ sky130_fd_sc_hd__a31o_1
X_25908_ _27572_/CLK _25908_/D vssd1 vssd1 vccd1 vccd1 _25908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17690_ _25916_/Q _17689_/X _17690_/S vssd1 vssd1 vccd1 vccd1 _17691_/A sky130_fd_sc_hd__mux2_1
X_26888_ _22414_/X _26888_/D vssd1 vssd1 vccd1 vccd1 _26888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16641_ _16641_/A vssd1 vssd1 vccd1 vccd1 _16877_/A sky130_fd_sc_hd__clkbuf_2
X_25839_ _26038_/CLK _25839_/D vssd1 vssd1 vccd1 vccd1 _25839_/Q sky130_fd_sc_hd__dfxtp_1
X_13853_ _15335_/A _14149_/B vssd1 vssd1 vccd1 vccd1 _13872_/A sky130_fd_sc_hd__or2_2
XFILLER_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19360_ _19469_/A vssd1 vssd1 vccd1 vccd1 _19360_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16572_ _16798_/B _16572_/B vssd1 vssd1 vccd1 vccd1 _16572_/X sky130_fd_sc_hd__and2_1
X_13784_ _26867_/Q _13778_/X _13780_/X _13783_/Y vssd1 vssd1 vccd1 vccd1 _26867_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18311_ _18468_/A vssd1 vssd1 vccd1 vccd1 _18311_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15523_ _13166_/X _26214_/Q _15523_/S vssd1 vssd1 vccd1 vccd1 _15524_/A sky130_fd_sc_hd__mux2_1
X_27509_ _27711_/CLK _27509_/D vssd1 vssd1 vccd1 vccd1 _27509_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19291_ _19282_/X _19285_/X _19289_/X _19290_/X _19220_/X vssd1 vssd1 vccd1 vccd1
+ _19292_/C sky130_fd_sc_hd__a221o_1
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18242_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18242_/X sky130_fd_sc_hd__buf_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _26245_/Q _13385_/X _15462_/S vssd1 vssd1 vccd1 vccd1 _15455_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14405_ _14441_/A vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18173_ _26951_/Q _26919_/Q _26887_/Q _26855_/Q _18101_/X _18129_/X vssd1 vssd1 vccd1
+ vccd1 _18173_/X sky130_fd_sc_hd__mux4_2
X_15385_ _15385_/A vssd1 vssd1 vccd1 vccd1 _26276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17124_ _17385_/S vssd1 vssd1 vccd1 vccd1 _17173_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14336_ _26679_/Q _14322_/X _14329_/X _14335_/Y vssd1 vssd1 vccd1 vccd1 _26679_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_117_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14267_ _26705_/Q _14256_/X _14258_/X _14266_/Y vssd1 vssd1 vccd1 vccd1 _26705_/D
+ sky130_fd_sc_hd__a31o_1
X_17055_ _17029_/X _17055_/B vssd1 vssd1 vccd1 vccd1 _17055_/X sky130_fd_sc_hd__and2b_1
XFILLER_125_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13218_ _13218_/A vssd1 vssd1 vccd1 vccd1 _27038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16006_ _16112_/B vssd1 vssd1 vccd1 vccd1 _16244_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14198_ _26729_/Q _14186_/X _14194_/X _14197_/Y vssd1 vssd1 vccd1 vccd1 _26729_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _27350_/Q _13061_/A _13081_/A _27318_/Q _13148_/X vssd1 vssd1 vccd1 vccd1
+ _16252_/A sky130_fd_sc_hd__a221o_4
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17957_ _17888_/X _17954_/X _17956_/X _17894_/X vssd1 vssd1 vccd1 vccd1 _17957_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater303 _27663_/CLK vssd1 vssd1 vccd1 vccd1 _27659_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater314 _27703_/CLK vssd1 vssd1 vccd1 vccd1 _27705_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater325 _27250_/CLK vssd1 vssd1 vccd1 vccd1 _27633_/CLK sky130_fd_sc_hd__clkbuf_1
X_16908_ _16908_/A _16908_/B vssd1 vssd1 vccd1 vccd1 _16908_/Y sky130_fd_sc_hd__nor2_1
Xrepeater336 _27782_/CLK vssd1 vssd1 vccd1 vccd1 _27781_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater347 _27645_/CLK vssd1 vssd1 vccd1 vccd1 _27753_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17888_ _18479_/A vssd1 vssd1 vccd1 vccd1 _17888_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater358 _27348_/CLK vssd1 vssd1 vccd1 vccd1 _27542_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater369 _27677_/CLK vssd1 vssd1 vccd1 vccd1 _27209_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19627_ _19621_/X _19622_/X _19623_/X _19624_/X _19625_/X _19626_/X vssd1 vssd1 vccd1
+ vccd1 _19628_/A sky130_fd_sc_hd__mux4_1
X_16839_ _16308_/A _16304_/A _16793_/A _16838_/Y vssd1 vssd1 vccd1 vccd1 _16839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19558_ _18801_/X _19553_/X _19555_/X _19557_/X _19312_/S vssd1 vssd1 vccd1 vccd1
+ _19567_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18509_ _18509_/A _18509_/B _18509_/C vssd1 vssd1 vccd1 vccd1 _18510_/A sky130_fd_sc_hd__and3_1
XFILLER_62_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ _19485_/X _19487_/X _19488_/X vssd1 vssd1 vccd1 vccd1 _19489_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21520_ _21520_/A vssd1 vssd1 vccd1 vccd1 _21520_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21451_ _21443_/X _21444_/X _21445_/X _21446_/X _21447_/X _21448_/X vssd1 vssd1 vccd1
+ vccd1 _21452_/A sky130_fd_sc_hd__mux4_1
XFILLER_193_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20402_ _20392_/X _20393_/X _20394_/X _20395_/X _20396_/X _20397_/X vssd1 vssd1 vccd1
+ vccd1 _20403_/A sky130_fd_sc_hd__mux4_1
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24170_ _24170_/A vssd1 vssd1 vccd1 vccd1 _27356_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_21382_ _21382_/A vssd1 vssd1 vccd1 vccd1 _21382_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23121_ _27102_/Q _17689_/X _23121_/S vssd1 vssd1 vccd1 vccd1 _23122_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_428 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20333_ _20333_/A vssd1 vssd1 vccd1 vccd1 _20333_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23052_ _23052_/A vssd1 vssd1 vccd1 vccd1 _27071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20264_ _20248_/X _20249_/X _20250_/X _20251_/X _20253_/X _20255_/X vssd1 vssd1 vccd1
+ vccd1 _20265_/A sky130_fd_sc_hd__mux4_1
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22003_ _22089_/A vssd1 vssd1 vccd1 vccd1 _22072_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20195_ _20195_/A vssd1 vssd1 vccd1 vccd1 _20195_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26811_ _22150_/X _26811_/D vssd1 vssd1 vccd1 vccd1 _26811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27791_ _27791_/CLK _27791_/D vssd1 vssd1 vccd1 vccd1 _27981_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_103_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26742_ _21906_/X _26742_/D vssd1 vssd1 vccd1 vccd1 _26742_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23954_ _24001_/A vssd1 vssd1 vccd1 vccd1 _23954_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22905_ _22888_/X _22890_/X _22892_/X _22894_/X _22895_/X _22896_/X vssd1 vssd1 vccd1
+ vccd1 _22906_/A sky130_fd_sc_hd__mux4_1
XFILLER_186_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26673_ _21662_/X _26673_/D vssd1 vssd1 vccd1 vccd1 _26673_/Q sky130_fd_sc_hd__dfxtp_1
X_23885_ _27079_/Q _27111_/Q _23892_/S vssd1 vssd1 vccd1 vccd1 _23885_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25624_ _25624_/A vssd1 vssd1 vccd1 vccd1 _27791_/D sky130_fd_sc_hd__clkbuf_1
X_22836_ _22836_/A vssd1 vssd1 vccd1 vccd1 _22836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25555_ _25547_/X _25552_/X _25553_/X _24920_/B _25554_/X vssd1 vssd1 vccd1 vccd1
+ _25555_/X sky130_fd_sc_hd__o311a_1
X_22767_ _22783_/A vssd1 vssd1 vccd1 vccd1 _22767_/X sky130_fd_sc_hd__clkbuf_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21718_ _21718_/A vssd1 vssd1 vccd1 vccd1 _21718_/X sky130_fd_sc_hd__clkbuf_1
X_24506_ _24407_/A _24633_/C _24505_/X _19313_/A vssd1 vssd1 vccd1 vccd1 _27523_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25486_ _27698_/Q _25479_/X _25480_/X vssd1 vssd1 vccd1 vccd1 _25486_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22698_ _22698_/A vssd1 vssd1 vccd1 vccd1 _22698_/X sky130_fd_sc_hd__clkbuf_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27225_ _27225_/CLK _27225_/D vssd1 vssd1 vccd1 vccd1 _27225_/Q sky130_fd_sc_hd__dfxtp_1
X_21649_ _21649_/A vssd1 vssd1 vccd1 vccd1 _21649_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_184_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24437_ _27617_/Q _24445_/B vssd1 vssd1 vccd1 vccd1 _24438_/A sky130_fd_sc_hd__and2_1
XFILLER_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15170_ _15170_/A vssd1 vssd1 vccd1 vccd1 _26371_/D sky130_fd_sc_hd__clkbuf_1
X_27156_ _27852_/CLK _27156_/D vssd1 vssd1 vccd1 vccd1 _27156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24368_ _27566_/Q _24372_/B vssd1 vssd1 vccd1 vccd1 _24369_/A sky130_fd_sc_hd__and2_1
XFILLER_193_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_90 _18944_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _14386_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26107_ _19689_/X _26107_/D vssd1 vssd1 vccd1 vccd1 _26107_/Q sky130_fd_sc_hd__dfxtp_1
X_23319_ _27728_/Q _23315_/Y _27732_/Q _23284_/Y _23318_/X vssd1 vssd1 vccd1 vccd1
+ _23319_/X sky130_fd_sc_hd__o221a_1
XFILLER_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27087_ _27295_/CLK _27087_/D vssd1 vssd1 vccd1 vccd1 _27087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24299_ _16287_/X _16288_/Y _16289_/X _25618_/B vssd1 vssd1 vccd1 vccd1 _27429_/D
+ sky130_fd_sc_hd__a31oi_4
XFILLER_153_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _14524_/A vssd1 vssd1 vccd1 vccd1 _14408_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26038_ _26038_/CLK _26038_/D vssd1 vssd1 vccd1 vccd1 _26038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ _27797_/Q _13009_/B vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__and2_1
X_18860_ _26267_/Q _26235_/Q _26203_/Q _26171_/Q _18859_/X _18818_/X vssd1 vssd1 vccd1
+ vccd1 _18860_/X sky130_fd_sc_hd__mux4_1
X_17811_ _26682_/Q _26650_/Q _26618_/Q _26586_/Q _18387_/A _17810_/X vssd1 vssd1 vccd1
+ vccd1 _17814_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27950__436 vssd1 vssd1 vccd1 vccd1 _27950__436/HI _27950_/A sky130_fd_sc_hd__conb_1
X_18791_ _26938_/Q _26906_/Q _26874_/Q _26842_/Q _18788_/X _18790_/X vssd1 vssd1 vccd1
+ vccd1 _18791_/X sky130_fd_sc_hd__mux4_2
XFILLER_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27989_ _27989_/A _15893_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_17742_ _25932_/Q _17740_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17743_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14954_ _14954_/A vssd1 vssd1 vccd1 vccd1 _26459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13905_ _26824_/Q _13893_/X _13899_/X _13904_/Y vssd1 vssd1 vccd1 vccd1 _26824_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_36_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17673_ _27408_/Q vssd1 vssd1 vccd1 vccd1 _17673_/X sky130_fd_sc_hd__clkbuf_2
X_14885_ _14885_/A _15783_/B vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__or2_2
XFILLER_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19412_ _19412_/A vssd1 vssd1 vccd1 vccd1 _19412_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16624_ _16621_/X _16804_/B _16804_/A vssd1 vssd1 vccd1 vccd1 _16624_/X sky130_fd_sc_hd__o21ba_1
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13836_ _13928_/A _13838_/B vssd1 vssd1 vccd1 vccd1 _13836_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_565 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19343_/A vssd1 vssd1 vccd1 vccd1 _19343_/X sky130_fd_sc_hd__buf_2
X_16555_ _16700_/A _16514_/X _16542_/X _16554_/X vssd1 vssd1 vccd1 vccd1 _16888_/A
+ sky130_fd_sc_hd__a31o_1
X_13767_ _26873_/Q _13761_/X _13764_/X _13766_/Y vssd1 vssd1 vccd1 vccd1 _26873_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_16_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ _13122_/X _26222_/Q _15512_/S vssd1 vssd1 vccd1 vccd1 _15507_/A sky130_fd_sc_hd__mux2_1
X_19274_ _26700_/Q _26668_/Q _26636_/Q _26604_/Q _19179_/X _19227_/X vssd1 vssd1 vccd1
+ vccd1 _19274_/X sky130_fd_sc_hd__mux4_2
XFILLER_149_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16486_ _16486_/A _16697_/A vssd1 vssd1 vccd1 vccd1 _16489_/C sky130_fd_sc_hd__nand2_1
X_13698_ _13878_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18225_ _26825_/Q _26793_/Q _26761_/Q _26729_/Q _18085_/X _17913_/X vssd1 vssd1 vccd1
+ vccd1 _18225_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15437_ _15437_/A vssd1 vssd1 vccd1 vccd1 _26253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18156_ _18156_/A vssd1 vssd1 vccd1 vccd1 _18156_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15368_ _14756_/X _26283_/Q _15368_/S vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17107_ _17094_/X _17107_/B vssd1 vssd1 vccd1 vccd1 _17107_/X sky130_fd_sc_hd__and2b_1
X_14319_ _26685_/Q _14310_/X _14311_/X _14318_/Y vssd1 vssd1 vccd1 vccd1 _26685_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18087_ _18009_/X _18086_/X _18014_/X vssd1 vssd1 vccd1 vccd1 _18087_/X sky130_fd_sc_hd__o21a_1
X_15299_ _15299_/A vssd1 vssd1 vccd1 vccd1 _26314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17038_ _27197_/Q _17037_/X _17067_/S vssd1 vssd1 vccd1 vccd1 _17039_/A sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater100 _27787_/CLK vssd1 vssd1 vccd1 vccd1 _27219_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _18989_/A _18989_/B _18989_/C vssd1 vssd1 vccd1 vccd1 _18990_/A sky130_fd_sc_hd__and3_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater111 _27122_/CLK vssd1 vssd1 vccd1 vccd1 _27126_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater122 _27788_/CLK vssd1 vssd1 vccd1 vccd1 _27675_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater133 _27845_/CLK vssd1 vssd1 vccd1 vccd1 _27844_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater144 _27211_/CLK vssd1 vssd1 vccd1 vccd1 _27127_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater155 _27407_/CLK vssd1 vssd1 vccd1 vccd1 _27383_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater166 _27789_/CLK vssd1 vssd1 vccd1 vccd1 _27792_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater177 _27110_/CLK vssd1 vssd1 vccd1 vccd1 _27111_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
X_20951_ _20937_/X _20938_/X _20939_/X _20940_/X _20941_/X _20942_/X vssd1 vssd1 vccd1
+ vccd1 _20952_/A sky130_fd_sc_hd__mux4_1
XFILLER_22_1169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xrepeater188 _26014_/CLK vssd1 vssd1 vccd1 vccd1 _27415_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater199 _27141_/CLK vssd1 vssd1 vccd1 vccd1 _25989_/CLK sky130_fd_sc_hd__clkbuf_1
X_23670_ _27761_/Q _27241_/Q _23672_/S vssd1 vssd1 vccd1 vccd1 _23671_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20882_ _20882_/A vssd1 vssd1 vccd1 vccd1 _20882_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22621_ _22609_/X _22610_/X _22611_/X _22612_/X _22615_/X _22618_/X vssd1 vssd1 vccd1
+ vccd1 _22622_/A sky130_fd_sc_hd__mux4_1
XFILLER_81_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25340_ _25347_/A _27516_/Q vssd1 vssd1 vccd1 vccd1 _25342_/A sky130_fd_sc_hd__nor2_1
X_22552_ _22552_/A vssd1 vssd1 vccd1 vccd1 _22552_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_924 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21503_ _21494_/X _21496_/X _21498_/X _21500_/X _21501_/X _21502_/X vssd1 vssd1 vccd1
+ vccd1 _21504_/A sky130_fd_sc_hd__mux4_1
X_25271_ _25272_/A _25272_/B _25272_/C vssd1 vssd1 vccd1 vccd1 _25273_/A sky130_fd_sc_hd__a21oi_2
X_22483_ _22471_/X _22472_/X _22473_/X _22474_/X _22475_/X _22476_/X vssd1 vssd1 vccd1
+ vccd1 _22484_/A sky130_fd_sc_hd__mux4_1
X_27010_ _22844_/X _27010_/D vssd1 vssd1 vccd1 vccd1 _27010_/Q sky130_fd_sc_hd__dfxtp_1
X_24222_ _25618_/A _24222_/B vssd1 vssd1 vccd1 vccd1 _27381_/D sky130_fd_sc_hd__nor2_1
X_21434_ _21434_/A vssd1 vssd1 vccd1 vccd1 _21434_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24153_ _24175_/A vssd1 vssd1 vccd1 vccd1 _24162_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21365_ _21357_/X _21358_/X _21359_/X _21360_/X _21361_/X _21362_/X vssd1 vssd1 vccd1
+ vccd1 _21366_/A sky130_fd_sc_hd__mux4_1
XFILLER_190_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23104_ _23104_/A vssd1 vssd1 vccd1 vccd1 _27095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20316_ _20302_/X _20303_/X _20304_/X _20305_/X _20306_/X _20307_/X vssd1 vssd1 vccd1
+ vccd1 _20317_/A sky130_fd_sc_hd__mux4_1
X_24084_ _27391_/Q _24084_/B vssd1 vssd1 vccd1 vccd1 _24085_/A sky130_fd_sc_hd__and2_1
X_21296_ _21296_/A vssd1 vssd1 vccd1 vccd1 _21296_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23035_ _23035_/A _27382_/Q _23035_/C _23035_/D vssd1 vssd1 vccd1 vccd1 _23109_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_192_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20247_ _20247_/A vssd1 vssd1 vccd1 vccd1 _20247_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27843_ _27845_/CLK _27843_/D vssd1 vssd1 vccd1 vccd1 _27843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20178_ _20162_/X _20163_/X _20164_/X _20165_/X _20167_/X _20169_/X vssd1 vssd1 vccd1
+ vccd1 _20179_/A sky130_fd_sc_hd__mux4_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27774_ _27774_/CLK _27774_/D vssd1 vssd1 vccd1 vccd1 _27774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24986_ _27067_/Q _27099_/Q _25004_/S vssd1 vssd1 vccd1 vccd1 _24986_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26725_ _21854_/X _26725_/D vssd1 vssd1 vccd1 vccd1 _26725_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23937_ _25931_/Q _25997_/Q _25830_/Q _26029_/Q _23899_/X _23929_/X vssd1 vssd1 vccd1
+ vccd1 _23937_/X sky130_fd_sc_hd__mux4_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26656_ _21608_/X _26656_/D vssd1 vssd1 vccd1 vccd1 _26656_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _26569_/Q _14658_/X _14666_/X _14669_/Y vssd1 vssd1 vccd1 vccd1 _26569_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23868_ _23866_/X _23867_/X _23891_/S vssd1 vssd1 vccd1 vccd1 _23868_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _13891_/A _13621_/B vssd1 vssd1 vccd1 vccd1 _13621_/Y sky130_fd_sc_hd__nor2_1
X_25607_ _25517_/A _25582_/X _25583_/X _24967_/B _25584_/X vssd1 vssd1 vccd1 vccd1
+ _25607_/X sky130_fd_sc_hd__o311a_1
XFILLER_60_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22819_ _22802_/X _22804_/X _22806_/X _22808_/X _22809_/X _22810_/X vssd1 vssd1 vccd1
+ vccd1 _22820_/A sky130_fd_sc_hd__mux4_1
X_26587_ _21368_/X _26587_/D vssd1 vssd1 vccd1 vccd1 _26587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23799_ _23740_/X _23797_/X _23798_/X _23768_/X vssd1 vssd1 vccd1 vccd1 _27275_/D
+ sky130_fd_sc_hd__o211a_1
X_16340_ _14810_/A _16501_/A _16374_/A _25944_/Q _16339_/X vssd1 vssd1 vccd1 vccd1
+ _16759_/B sky130_fd_sc_hd__a221o_2
X_13552_ _26945_/Q _13535_/X _13528_/X _13551_/Y vssd1 vssd1 vccd1 vccd1 _26945_/D
+ sky130_fd_sc_hd__a31o_1
X_25538_ _24778_/A _25534_/X _25535_/Y _25537_/X _25527_/X vssd1 vssd1 vccd1 vccd1
+ _27770_/D sky130_fd_sc_hd__a221oi_1
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16271_ _16271_/A _16276_/B _16296_/B vssd1 vssd1 vccd1 vccd1 _16271_/X sky130_fd_sc_hd__and3_1
X_13483_ _27356_/Q _13062_/A _13082_/A _27324_/Q _13114_/X vssd1 vssd1 vccd1 vccd1
+ _16289_/A sky130_fd_sc_hd__a221oi_4
XFILLER_201_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25469_ _27695_/Q _25448_/X _25449_/X vssd1 vssd1 vccd1 vccd1 _25469_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18010_ _18177_/A vssd1 vssd1 vccd1 vccd1 _18011_/A sky130_fd_sc_hd__buf_6
XFILLER_139_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15222_ _15222_/A vssd1 vssd1 vccd1 vccd1 _26348_/D sky130_fd_sc_hd__clkbuf_1
X_27208_ _27208_/CLK _27208_/D vssd1 vssd1 vccd1 vccd1 _27208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1045 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27139_ _27140_/CLK _27139_/D vssd1 vssd1 vccd1 vccd1 _27139_/Q sky130_fd_sc_hd__dfxtp_1
X_15153_ _15175_/A vssd1 vssd1 vccd1 vccd1 _15162_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_181_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14104_ _14157_/A vssd1 vssd1 vccd1 vccd1 _14104_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15084_ _14763_/X _26409_/Q _15090_/S vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19961_ _19977_/A vssd1 vssd1 vccd1 vccd1 _19961_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14035_ _14507_/A vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18912_ _18929_/A vssd1 vssd1 vccd1 vccd1 _24403_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19892_ _19882_/X _19883_/X _19884_/X _19885_/X _19886_/X _19887_/X vssd1 vssd1 vccd1
+ vccd1 _19893_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18843_ _18843_/A vssd1 vssd1 vccd1 vccd1 _26042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18774_ _19296_/S vssd1 vssd1 vccd1 vccd1 _19553_/S sky130_fd_sc_hd__buf_4
XFILLER_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15986_ _15988_/A vssd1 vssd1 vccd1 vccd1 _15986_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _17757_/A vssd1 vssd1 vccd1 vccd1 _17738_/S sky130_fd_sc_hd__buf_2
XFILLER_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14937_ _14937_/A vssd1 vssd1 vccd1 vccd1 _26467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17656_ _17501_/X _25899_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _17657_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14868_ _26497_/Q _13398_/X _14868_/S vssd1 vssd1 vccd1 vccd1 _14869_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16607_ _16481_/A _16606_/Y _16686_/A _16450_/Y vssd1 vssd1 vccd1 vccd1 _16692_/A
+ sky130_fd_sc_hd__a211oi_1
X_13819_ _13844_/A vssd1 vssd1 vccd1 vccd1 _13819_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17587_ _17504_/X _25868_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17588_/A sky130_fd_sc_hd__mux2_1
X_14799_ _14798_/X _26526_/Q _14805_/S vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19326_ _19460_/A vssd1 vssd1 vccd1 vccd1 _19326_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16538_ _16822_/A vssd1 vssd1 vccd1 vccd1 _16616_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19257_ _19254_/X _19256_/X _19346_/S vssd1 vssd1 vccd1 vccd1 _19257_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16469_ _16611_/B _16469_/B vssd1 vssd1 vccd1 vccd1 _16469_/X sky130_fd_sc_hd__and2_1
X_18208_ _18208_/A _18207_/X vssd1 vssd1 vccd1 vccd1 _18208_/X sky130_fd_sc_hd__or2b_1
XFILLER_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19188_ _19482_/A vssd1 vssd1 vccd1 vccd1 _19188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18139_ _26277_/Q _26245_/Q _26213_/Q _26181_/Q _18044_/X _18068_/X vssd1 vssd1 vccd1
+ vccd1 _18139_/X sky130_fd_sc_hd__mux4_2
XFILLER_89_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21150_ _21214_/A vssd1 vssd1 vccd1 vccd1 _21150_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20101_ _20165_/A vssd1 vssd1 vccd1 vccd1 _20101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21081_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21081_/X sky130_fd_sc_hd__clkbuf_2
X_20032_ _20064_/A vssd1 vssd1 vccd1 vccd1 _20032_/X sky130_fd_sc_hd__clkbuf_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24840_ _27644_/Q _24834_/X _24838_/Y _24839_/X vssd1 vssd1 vccd1 vccd1 _27644_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21983_ _21999_/A vssd1 vssd1 vccd1 vccd1 _21983_/X sky130_fd_sc_hd__clkbuf_1
X_24771_ _24771_/A vssd1 vssd1 vccd1 vccd1 _24771_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26510_ _21100_/X _26510_/D vssd1 vssd1 vccd1 vccd1 _26510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ _20934_/A vssd1 vssd1 vccd1 vccd1 _20934_/X sky130_fd_sc_hd__clkbuf_1
X_23722_ _27825_/Q _25358_/A vssd1 vssd1 vccd1 vccd1 _24186_/A sky130_fd_sc_hd__nor2_2
XFILLER_82_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27490_ _27534_/CLK _27490_/D vssd1 vssd1 vccd1 vccd1 _27490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26441_ _20857_/X _26441_/D vssd1 vssd1 vccd1 vccd1 _26441_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20865_/X sky130_fd_sc_hd__clkbuf_1
X_23653_ _25976_/Q _27233_/Q _23661_/S vssd1 vssd1 vccd1 vccd1 _23654_/A sky130_fd_sc_hd__mux2_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22604_ _22604_/A vssd1 vssd1 vccd1 vccd1 _22604_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23584_ _27774_/Q vssd1 vssd1 vccd1 vccd1 _24925_/B sky130_fd_sc_hd__buf_4
X_26372_ _20611_/X _26372_/D vssd1 vssd1 vccd1 vccd1 _26372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20796_ _20796_/A vssd1 vssd1 vccd1 vccd1 _22543_/A sky130_fd_sc_hd__buf_6
XFILLER_167_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22535_ _22519_/X _22520_/X _22521_/X _22522_/X _22524_/X _22526_/X vssd1 vssd1 vccd1
+ vccd1 _22536_/A sky130_fd_sc_hd__mux4_1
X_25323_ _25323_/A _27514_/Q vssd1 vssd1 vccd1 vccd1 _25325_/A sky130_fd_sc_hd__xor2_1
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22466_ _22466_/A vssd1 vssd1 vccd1 vccd1 _22466_/X sky130_fd_sc_hd__clkbuf_1
X_25254_ _25297_/A vssd1 vssd1 vccd1 vccd1 _25254_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21417_ _21408_/X _21410_/X _21412_/X _21414_/X _21415_/X _21416_/X vssd1 vssd1 vccd1
+ vccd1 _21418_/A sky130_fd_sc_hd__mux4_1
X_24205_ _24217_/A vssd1 vssd1 vccd1 vccd1 _24210_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25185_ _25309_/A vssd1 vssd1 vccd1 vccd1 _25221_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22397_ _22385_/X _22386_/X _22387_/X _22388_/X _22389_/X _22390_/X vssd1 vssd1 vccd1
+ vccd1 _22398_/A sky130_fd_sc_hd__mux4_1
XFILLER_136_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24136_ _27446_/Q _24140_/B vssd1 vssd1 vccd1 vccd1 _24137_/A sky130_fd_sc_hd__and2_1
X_21348_ _21348_/A vssd1 vssd1 vccd1 vccd1 _21348_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24067_ _24067_/A vssd1 vssd1 vccd1 vccd1 _27310_/D sky130_fd_sc_hd__clkbuf_1
X_21279_ _21269_/X _21270_/X _21271_/X _21272_/X _21273_/X _21274_/X vssd1 vssd1 vccd1
+ vccd1 _21280_/A sky130_fd_sc_hd__mux4_1
X_23018_ _23018_/A vssd1 vssd1 vccd1 vccd1 _23018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27826_ _27826_/CLK _27826_/D vssd1 vssd1 vccd1 vccd1 _27826_/Q sky130_fd_sc_hd__dfxtp_1
X_15840_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15849_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15771_/A _15771_/B vssd1 vssd1 vccd1 vccd1 _15771_/Y sky130_fd_sc_hd__nor2_1
X_27757_ _27758_/CLK _27757_/D vssd1 vssd1 vccd1 vccd1 _27757_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _27806_/Q _12987_/B vssd1 vssd1 vccd1 vccd1 _12984_/A sky130_fd_sc_hd__and2_1
X_24969_ _24969_/A _24969_/B vssd1 vssd1 vccd1 vccd1 _24970_/B sky130_fd_sc_hd__xnor2_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17510_ _17510_/A vssd1 vssd1 vccd1 vccd1 _25837_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26708_ _21790_/X _26708_/D vssd1 vssd1 vccd1 vccd1 _26708_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14722_ _14721_/X _26550_/Q _14725_/S vssd1 vssd1 vccd1 vccd1 _14723_/A sky130_fd_sc_hd__mux2_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ _18480_/X _18484_/X _18488_/X _18443_/X _18489_/X vssd1 vssd1 vccd1 vccd1
+ _18491_/C sky130_fd_sc_hd__a221o_1
XFILLER_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27688_ _27753_/CLK _27688_/D vssd1 vssd1 vccd1 vccd1 _27688_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17524_/S vssd1 vssd1 vccd1 vccd1 _17454_/S sky130_fd_sc_hd__clkbuf_2
X_26639_ _21544_/X _26639_/D vssd1 vssd1 vccd1 vccd1 _26639_/Q sky130_fd_sc_hd__dfxtp_1
X_14653_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14653_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13604_ _13874_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13604_/Y sky130_fd_sc_hd__nor2_1
X_17372_ _25841_/Q _26040_/Q _17382_/S vssd1 vssd1 vccd1 vccd1 _17372_/X sky130_fd_sc_hd__mux2_1
X_14584_ _15745_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14584_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19111_ _19407_/A vssd1 vssd1 vccd1 vccd1 _19111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16323_ _17410_/A _16490_/B vssd1 vssd1 vccd1 vccd1 _16323_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ _13558_/A vssd1 vssd1 vccd1 vccd1 _13535_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19042_ _26690_/Q _26658_/Q _26626_/Q _26594_/Q _19015_/X _18939_/X vssd1 vssd1 vccd1
+ vccd1 _19042_/X sky130_fd_sc_hd__mux4_2
XFILLER_146_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16254_ _24290_/A _27534_/Q _16254_/S vssd1 vssd1 vccd1 vccd1 _16453_/A sky130_fd_sc_hd__mux2_1
X_13466_ _16298_/A vssd1 vssd1 vccd1 vccd1 _13876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_185_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15205_ _15205_/A vssd1 vssd1 vccd1 vccd1 _26356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16185_ _26042_/Q _16215_/B _16221_/C _16184_/X vssd1 vssd1 vccd1 vccd1 _16185_/X
+ sky130_fd_sc_hd__a31o_1
X_13397_ _13397_/A vssd1 vssd1 vccd1 vccd1 _26978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15136_ _26386_/Q _13344_/X _15140_/S vssd1 vssd1 vccd1 vccd1 _15137_/A sky130_fd_sc_hd__mux2_1
X_27956__442 vssd1 vssd1 vccd1 vccd1 _27956__442/HI _27956_/A sky130_fd_sc_hd__conb_1
XFILLER_153_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15067_ _15067_/A vssd1 vssd1 vccd1 vccd1 _26417_/D sky130_fd_sc_hd__clkbuf_1
X_19944_ _19976_/A vssd1 vssd1 vccd1 vccd1 _19944_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _26790_/Q _14005_/X _14001_/X _14017_/Y vssd1 vssd1 vccd1 vccd1 _26790_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19875_ _19875_/A vssd1 vssd1 vccd1 vccd1 _19875_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18826_ _19399_/A vssd1 vssd1 vccd1 vccd1 _18826_/X sky130_fd_sc_hd__buf_4
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18757_ _26039_/Q _17769_/X _18757_/S vssd1 vssd1 vccd1 vccd1 _18758_/A sky130_fd_sc_hd__mux2_1
X_15969_ _15973_/A vssd1 vssd1 vccd1 vccd1 _15969_/Y sky130_fd_sc_hd__inv_2
X_17708_ _27418_/Q vssd1 vssd1 vccd1 vccd1 _17708_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18688_ _18688_/A vssd1 vssd1 vccd1 vccd1 _26008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ _17476_/X _25891_/Q _17645_/S vssd1 vssd1 vccd1 vccd1 _17640_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20650_ _20636_/X _20637_/X _20638_/X _20639_/X _20640_/X _20641_/X vssd1 vssd1 vccd1
+ vccd1 _20651_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _19307_/X _19308_/X _19492_/A vssd1 vssd1 vccd1 vccd1 _19309_/X sky130_fd_sc_hd__mux2_2
XFILLER_56_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20581_ _20581_/A vssd1 vssd1 vccd1 vccd1 _20581_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22320_ _22336_/A vssd1 vssd1 vccd1 vccd1 _22320_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22251_ _22245_/X _22246_/X _22247_/X _22248_/X _22249_/X _22250_/X vssd1 vssd1 vccd1
+ vccd1 _22252_/A sky130_fd_sc_hd__mux4_1
XFILLER_118_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21202_ _21202_/A vssd1 vssd1 vccd1 vccd1 _21202_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22182_ _22250_/A vssd1 vssd1 vccd1 vccd1 _22182_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21133_ _21125_/X _21126_/X _21127_/X _21128_/X _21130_/X _21132_/X vssd1 vssd1 vccd1
+ vccd1 _21134_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26990_ _22774_/X _26990_/D vssd1 vssd1 vccd1 vccd1 _26990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25941_ _25941_/CLK _25941_/D vssd1 vssd1 vccd1 vccd1 _25941_/Q sky130_fd_sc_hd__dfxtp_1
X_21064_ _21128_/A vssd1 vssd1 vccd1 vccd1 _21064_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20015_ _20079_/A vssd1 vssd1 vccd1 vccd1 _20015_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25872_ _27854_/CLK _25872_/D vssd1 vssd1 vccd1 vccd1 _25872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27611_ _27611_/CLK _27611_/D vssd1 vssd1 vccd1 vccd1 _27611_/Q sky130_fd_sc_hd__dfxtp_1
X_24823_ _24823_/A _25601_/B vssd1 vssd1 vccd1 vccd1 _24823_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27542_ _27542_/CLK _27542_/D vssd1 vssd1 vccd1 vccd1 _27542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24754_ _24754_/A _24759_/B vssd1 vssd1 vccd1 vccd1 _24754_/Y sky130_fd_sc_hd__nand2_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21966_ _21998_/A vssd1 vssd1 vccd1 vccd1 _21966_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23705_ _25580_/A _27257_/Q _23705_/S vssd1 vssd1 vccd1 vccd1 _23706_/A sky130_fd_sc_hd__mux2_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27473_ _27473_/CLK _27473_/D vssd1 vssd1 vccd1 vccd1 _27473_/Q sky130_fd_sc_hd__dfxtp_1
X_20917_ _20905_/X _20906_/X _20907_/X _20908_/X _20909_/X _20910_/X vssd1 vssd1 vccd1
+ vccd1 _20918_/A sky130_fd_sc_hd__mux4_1
X_21897_ _21913_/A vssd1 vssd1 vccd1 vccd1 _21897_/X sky130_fd_sc_hd__clkbuf_1
X_24685_ _27176_/Q _24685_/B vssd1 vssd1 vccd1 vccd1 _24685_/X sky130_fd_sc_hd__or2_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26424_ _20787_/X _26424_/D vssd1 vssd1 vccd1 vccd1 _26424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20848_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20848_/X sky130_fd_sc_hd__clkbuf_1
X_23636_ _27230_/Q vssd1 vssd1 vccd1 vccd1 _25035_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26355_ _20557_/X _26355_/D vssd1 vssd1 vccd1 vccd1 _26355_/Q sky130_fd_sc_hd__dfxtp_1
X_23567_ _27769_/Q _27211_/Q _23576_/S vssd1 vssd1 vccd1 vccd1 _23568_/B sky130_fd_sc_hd__mux2_1
X_20779_ _20779_/A vssd1 vssd1 vccd1 vccd1 _20779_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25306_ _25306_/A _25306_/B vssd1 vssd1 vccd1 vccd1 _25306_/Y sky130_fd_sc_hd__nand2_1
X_13320_ _15551_/A _15783_/A vssd1 vssd1 vccd1 vccd1 _13402_/A sky130_fd_sc_hd__nor2_2
X_22518_ _22518_/A vssd1 vssd1 vccd1 vccd1 _22518_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23498_ _25132_/A vssd1 vssd1 vccd1 vccd1 _23498_/X sky130_fd_sc_hd__clkbuf_2
X_26286_ _20311_/X _26286_/D vssd1 vssd1 vccd1 vccd1 _26286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22449_ _22433_/X _22434_/X _22435_/X _22436_/X _22438_/X _22440_/X vssd1 vssd1 vccd1
+ vccd1 _22450_/A sky130_fd_sc_hd__mux4_1
X_25237_ _25261_/A _25237_/B vssd1 vssd1 vccd1 vccd1 _25237_/Y sky130_fd_sc_hd__nand2_1
X_13251_ _13251_/A vssd1 vssd1 vccd1 vccd1 _27033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13182_ _27280_/Q _13201_/B vssd1 vssd1 vccd1 vccd1 _13182_/X sky130_fd_sc_hd__and2_2
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25168_ _27527_/Q _27495_/Q vssd1 vssd1 vccd1 vccd1 _25170_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24119_ _24119_/A vssd1 vssd1 vccd1 vccd1 _24128_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25099_ _27841_/Q _27145_/Q _25890_/Q _25858_/Q _24974_/X _24975_/X vssd1 vssd1 vccd1
+ vccd1 _25099_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _18238_/A vssd1 vssd1 vccd1 vccd1 _17990_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16941_ _27600_/Q vssd1 vssd1 vccd1 vccd1 _18945_/A sky130_fd_sc_hd__inv_2
XFILLER_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19660_ _19832_/A vssd1 vssd1 vccd1 vccd1 _19727_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16872_ _24215_/A _25617_/A _25616_/A _16872_/D vssd1 vssd1 vccd1 vccd1 _16873_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18611_ _27541_/Q _27520_/Q vssd1 vssd1 vccd1 vccd1 _18612_/B sky130_fd_sc_hd__or2_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27809_ _25684_/X _27809_/D vssd1 vssd1 vccd1 vccd1 _27809_/Q sky130_fd_sc_hd__dfxtp_1
X_15823_ _13156_/X _26088_/Q _15827_/S vssd1 vssd1 vccd1 vccd1 _15824_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19591_ _19639_/A vssd1 vssd1 vccd1 vccd1 _19591_/X sky130_fd_sc_hd__clkbuf_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18542_ _26551_/Q _26519_/Q _26487_/Q _27063_/Q _17846_/X _17848_/X vssd1 vssd1 vccd1
+ vccd1 _18542_/X sky130_fd_sc_hd__mux4_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15754_/A _15758_/B vssd1 vssd1 vccd1 vccd1 _15754_/Y sky130_fd_sc_hd__nor2_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ _12966_/A vssd1 vssd1 vccd1 vccd1 _27814_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _15779_/A _14707_/B vssd1 vssd1 vccd1 vccd1 _14705_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18473_ _26708_/Q _26676_/Q _26644_/Q _26612_/Q _18360_/X _18408_/X vssd1 vssd1 vccd1
+ vccd1 _18475_/A sky130_fd_sc_hd__mux4_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15685_ _13216_/X _26142_/Q _15689_/S vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__mux2_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _14438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_361 _25659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17424_ _17505_/A vssd1 vssd1 vccd1 vccd1 _17524_/S sky130_fd_sc_hd__buf_2
XANTENNA_372 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_383 _16298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14636_ _26582_/Q _14630_/X _14624_/X _14635_/Y vssd1 vssd1 vccd1 vccd1 _26582_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17355_ _27094_/Q _27126_/Q _17355_/S vssd1 vssd1 vccd1 vccd1 _17355_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14567_ _15728_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14567_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16306_ _16576_/A _16304_/A _16304_/Y _16603_/A vssd1 vssd1 vccd1 vccd1 _16308_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13518_ _26952_/Q _13510_/X _13505_/X _13517_/Y vssd1 vssd1 vccd1 vccd1 _26952_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_201_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17286_ _27217_/Q _17285_/X _17311_/S vssd1 vssd1 vccd1 vccd1 _17287_/A sky130_fd_sc_hd__mux2_1
X_14498_ _15756_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _14498_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ _19299_/A vssd1 vssd1 vccd1 vccd1 _19123_/A sky130_fd_sc_hd__clkbuf_1
X_16237_ _15992_/A _16233_/X _16234_/X _16235_/X _16236_/X vssd1 vssd1 vccd1 vccd1
+ _16406_/A sky130_fd_sc_hd__o41a_1
XFILLER_174_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13449_ _26966_/Q _13435_/X _13429_/X _13448_/Y vssd1 vssd1 vccd1 vccd1 _26966_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16168_ _16426_/A _16252_/B vssd1 vssd1 vccd1 vccd1 _16168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_177_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15119_ _15175_/A vssd1 vssd1 vccd1 vccd1 _15188_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16099_ _16099_/A _16536_/B vssd1 vssd1 vccd1 vccd1 _16099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19927_ _19991_/A vssd1 vssd1 vccd1 vccd1 _19927_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19858_ _19850_/X _19851_/X _19852_/X _19853_/X _19854_/X _19855_/X vssd1 vssd1 vccd1
+ vccd1 _19859_/A sky130_fd_sc_hd__mux4_1
XFILLER_110_551 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18809_ _19401_/A vssd1 vssd1 vccd1 vccd1 _18926_/A sky130_fd_sc_hd__buf_2
X_19789_ _19789_/A vssd1 vssd1 vccd1 vccd1 _19789_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21820_ _21820_/A vssd1 vssd1 vccd1 vccd1 _21820_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21751_ _21737_/X _21738_/X _21739_/X _21740_/X _21743_/X _21746_/X vssd1 vssd1 vccd1
+ vccd1 _21752_/A sky130_fd_sc_hd__mux4_1
XFILLER_184_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20702_ _20702_/A vssd1 vssd1 vccd1 vccd1 _20770_/A sky130_fd_sc_hd__buf_2
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21682_ _21682_/A vssd1 vssd1 vccd1 vccd1 _21682_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24470_ _27632_/Q _24478_/B vssd1 vssd1 vccd1 vccd1 _24471_/A sky130_fd_sc_hd__and2_1
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20633_ _20633_/A vssd1 vssd1 vccd1 vccd1 _20633_/X sky130_fd_sc_hd__clkbuf_1
X_23421_ _23624_/A vssd1 vssd1 vccd1 vccd1 _23421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23352_ _24754_/A _27241_/Q _27253_/Q _24786_/A _23351_/Y vssd1 vssd1 vccd1 vccd1
+ _23360_/B sky130_fd_sc_hd__o221a_1
XFILLER_20_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26140_ _19803_/X _26140_/D vssd1 vssd1 vccd1 vccd1 _26140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20564_ _20550_/X _20551_/X _20552_/X _20553_/X _20554_/X _20555_/X vssd1 vssd1 vccd1
+ vccd1 _20565_/A sky130_fd_sc_hd__mux4_1
XFILLER_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22303_ _22335_/A vssd1 vssd1 vccd1 vccd1 _22303_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26071_ _27332_/CLK _26071_/D vssd1 vssd1 vccd1 vccd1 _26071_/Q sky130_fd_sc_hd__dfxtp_1
X_23283_ _23280_/Y input41/X _27723_/Q _23281_/Y _23282_/X vssd1 vssd1 vccd1 vccd1
+ _23293_/A sky130_fd_sc_hd__a221o_1
X_20495_ _20495_/A vssd1 vssd1 vccd1 vccd1 _20495_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22234_ _22250_/A vssd1 vssd1 vccd1 vccd1 _22234_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25022_ _27071_/Q _27103_/Q _25047_/S vssd1 vssd1 vccd1 vccd1 _25022_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22165_ _22157_/X _22158_/X _22159_/X _22160_/X _22161_/X _22162_/X vssd1 vssd1 vccd1
+ vccd1 _22166_/A sky130_fd_sc_hd__mux4_1
XFILLER_133_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21116_ _21116_/A vssd1 vssd1 vccd1 vccd1 _21116_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22096_ _22096_/A vssd1 vssd1 vccd1 vccd1 _22096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26973_ _22712_/X _26973_/D vssd1 vssd1 vccd1 vccd1 _26973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25924_ _25989_/CLK _25924_/D vssd1 vssd1 vccd1 vccd1 _25924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21047_ _21039_/X _21040_/X _21041_/X _21042_/X _21044_/X _21046_/X vssd1 vssd1 vccd1
+ vccd1 _21048_/A sky130_fd_sc_hd__mux4_1
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25855_ _27142_/CLK _25855_/D vssd1 vssd1 vccd1 vccd1 _25855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24806_ _24806_/A _24815_/B vssd1 vssd1 vccd1 vccd1 _24806_/Y sky130_fd_sc_hd__nand2_1
X_25786_ _17495_/X _27848_/Q _25790_/S vssd1 vssd1 vccd1 vccd1 _25787_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22998_ _23030_/A vssd1 vssd1 vccd1 vccd1 _22998_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27525_ _27529_/CLK _27525_/D vssd1 vssd1 vccd1 vccd1 _27525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24737_ _24737_/A _24970_/A vssd1 vssd1 vccd1 vccd1 _24737_/Y sky130_fd_sc_hd__nand2_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21949_ _21997_/A vssd1 vssd1 vccd1 vccd1 _21949_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_816 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27456_ _27458_/CLK _27456_/D vssd1 vssd1 vccd1 vccd1 _27456_/Q sky130_fd_sc_hd__dfxtp_1
X_15470_ _15470_/A vssd1 vssd1 vccd1 vccd1 _26238_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24668_ _27585_/Q _24660_/X _24667_/X _24663_/X vssd1 vssd1 vccd1 vccd1 _27585_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14441_/A vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26407_ _20733_/X _26407_/D vssd1 vssd1 vccd1 vccd1 _26407_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23619_ _27783_/Q vssd1 vssd1 vccd1 vccd1 _24965_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27387_ _27388_/CLK _27387_/D vssd1 vssd1 vccd1 vccd1 _27387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24599_ _24599_/A vssd1 vssd1 vccd1 vccd1 _27559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17140_ _27205_/Q _17138_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17141_/A sky130_fd_sc_hd__mux2_1
X_14352_ _14365_/A vssd1 vssd1 vccd1 vccd1 _14352_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26338_ _20493_/X _26338_/D vssd1 vssd1 vccd1 vccd1 _26338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13303_ _13303_/A vssd1 vssd1 vccd1 vccd1 _27009_/D sky130_fd_sc_hd__clkbuf_1
X_17071_ _25917_/Q _25983_/Q _17071_/S vssd1 vssd1 vccd1 vccd1 _17072_/B sky130_fd_sc_hd__mux2_1
X_14283_ _14296_/A vssd1 vssd1 vccd1 vccd1 _14283_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26269_ _20247_/X _26269_/D vssd1 vssd1 vccd1 vccd1 _26269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1058 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_28008_ _28008_/A _15858_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
X_16022_ _16205_/A vssd1 vssd1 vccd1 vccd1 _16197_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13234_ _14807_/A vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ _27347_/Q _13017_/A _13025_/A _27315_/Q _13164_/X vssd1 vssd1 vccd1 vccd1
+ _16240_/A sky130_fd_sc_hd__a221o_4
XFILLER_156_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17973_ _27798_/Q _26559_/Q _26431_/Q _26111_/Q _17920_/X _17949_/X vssd1 vssd1 vccd1
+ vccd1 _17973_/X sky130_fd_sc_hd__mux4_2
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13096_ _13096_/A vssd1 vssd1 vccd1 vccd1 _27059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19712_ _19728_/A vssd1 vssd1 vccd1 vccd1 _19712_/X sky130_fd_sc_hd__clkbuf_1
X_16924_ input2/X _27858_/Q vssd1 vssd1 vccd1 vccd1 _25358_/A sky130_fd_sc_hd__or2_4
XFILLER_46_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19643_ _25725_/A vssd1 vssd1 vccd1 vccd1 _19714_/A sky130_fd_sc_hd__buf_2
X_16855_ _16764_/A _16395_/A _16854_/X vssd1 vssd1 vccd1 vccd1 _16855_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15806_ _15806_/A vssd1 vssd1 vccd1 vccd1 _26096_/D sky130_fd_sc_hd__clkbuf_1
X_19574_ _19639_/A vssd1 vssd1 vccd1 vccd1 _19574_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16786_ _16786_/A _16786_/B _16722_/A vssd1 vssd1 vccd1 vccd1 _16786_/X sky130_fd_sc_hd__or3b_1
X_13998_ _14471_/A vssd1 vssd1 vccd1 vccd1 _14369_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18525_ _26294_/Q _26262_/Q _26230_/Q _26198_/Q _17801_/X _17805_/X vssd1 vssd1 vccd1
+ vccd1 _18525_/X sky130_fd_sc_hd__mux4_1
X_15737_ _26124_/Q _15734_/X _15727_/X _15736_/Y vssd1 vssd1 vccd1 vccd1 _26124_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12949_ _12949_/A vssd1 vssd1 vccd1 vccd1 _27821_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18456_ _26163_/Q _26099_/Q _27027_/Q _26995_/Q _18455_/X _18387_/X vssd1 vssd1 vccd1
+ vccd1 _18457_/A sky130_fd_sc_hd__mux4_2
X_15668_ _15668_/A vssd1 vssd1 vccd1 vccd1 _26150_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _16536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_191 _16451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17407_ _17407_/A vssd1 vssd1 vccd1 vccd1 _17407_/Y sky130_fd_sc_hd__clkinv_8
X_14619_ _26587_/Q _14615_/X _14542_/B _14618_/Y vssd1 vssd1 vccd1 vccd1 _26587_/D
+ sky130_fd_sc_hd__a31o_1
X_18387_ _18387_/A vssd1 vssd1 vccd1 vccd1 _18387_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15599_ _15599_/A vssd1 vssd1 vccd1 vccd1 _26181_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17338_ _17338_/A vssd1 vssd1 vccd1 vccd1 _17338_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17269_ _25832_/Q _26031_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17269_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19008_ _26528_/Q _26496_/Q _26464_/Q _27040_/Q _18984_/X _18863_/X vssd1 vssd1 vccd1
+ vccd1 _19008_/X sky130_fd_sc_hd__mux4_1
X_20280_ _20267_/X _20269_/X _20271_/X _20273_/X _20274_/X _20275_/X vssd1 vssd1 vccd1
+ vccd1 _20281_/A sky130_fd_sc_hd__mux4_1
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23970_ _23968_/X _23969_/X _23985_/S vssd1 vssd1 vccd1 vccd1 _23970_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22921_ _22907_/X _22908_/X _22909_/X _22910_/X _22911_/X _22912_/X vssd1 vssd1 vccd1
+ vccd1 _22922_/A sky130_fd_sc_hd__mux4_1
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25640_ _25709_/A vssd1 vssd1 vccd1 vccd1 _25640_/X sky130_fd_sc_hd__clkbuf_2
X_22852_ _22852_/A vssd1 vssd1 vccd1 vccd1 _22852_/X sky130_fd_sc_hd__clkbuf_1
X_21803_ _21793_/X _21794_/X _21795_/X _21796_/X _21797_/X _21798_/X vssd1 vssd1 vccd1
+ vccd1 _21804_/A sky130_fd_sc_hd__mux4_1
X_25571_ _24792_/A _25564_/X _25567_/X _25570_/Y _25557_/X vssd1 vssd1 vccd1 vccd1
+ _27775_/D sky130_fd_sc_hd__a221oi_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22783_ _22783_/A vssd1 vssd1 vccd1 vccd1 _22783_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27310_ _27311_/CLK _27310_/D vssd1 vssd1 vccd1 vccd1 _27310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24522_ _24522_/A _24631_/B vssd1 vssd1 vccd1 vccd1 _24522_/Y sky130_fd_sc_hd__nor2_1
X_21734_ _21734_/A vssd1 vssd1 vccd1 vccd1 _21734_/X sky130_fd_sc_hd__clkbuf_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27241_ _27258_/CLK _27241_/D vssd1 vssd1 vccd1 vccd1 _27241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24453_ _24453_/A vssd1 vssd1 vccd1 vccd1 _27503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21665_ _22537_/A vssd1 vssd1 vccd1 vccd1 _22015_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23404_ _27759_/Q vssd1 vssd1 vccd1 vccd1 _24848_/A sky130_fd_sc_hd__buf_2
XFILLER_184_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20616_ _20702_/A vssd1 vssd1 vccd1 vccd1 _20684_/A sky130_fd_sc_hd__clkbuf_2
X_27172_ _27172_/CLK _27172_/D vssd1 vssd1 vccd1 vccd1 _27172_/Q sky130_fd_sc_hd__dfxtp_1
X_21596_ _21596_/A vssd1 vssd1 vccd1 vccd1 _21596_/X sky130_fd_sc_hd__clkbuf_1
X_24384_ _24384_/A _24384_/B vssd1 vssd1 vccd1 vccd1 _27473_/D sky130_fd_sc_hd__nor2_1
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26123_ _19741_/X _26123_/D vssd1 vssd1 vccd1 vccd1 _26123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23335_ _27764_/Q vssd1 vssd1 vccd1 vccd1 _24763_/A sky130_fd_sc_hd__clkinv_2
X_20547_ _20547_/A vssd1 vssd1 vccd1 vccd1 _20547_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26054_ _26057_/CLK _26054_/D vssd1 vssd1 vccd1 vccd1 _26054_/Q sky130_fd_sc_hd__dfxtp_1
X_20478_ _20464_/X _20465_/X _20466_/X _20467_/X _20468_/X _20469_/X vssd1 vssd1 vccd1
+ vccd1 _20479_/A sky130_fd_sc_hd__mux4_1
X_23266_ _27743_/Q vssd1 vssd1 vccd1 vccd1 _23266_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25005_ _25003_/X _25004_/X _25031_/S vssd1 vssd1 vccd1 vccd1 _25005_/X sky130_fd_sc_hd__mux2_1
X_22217_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22217_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23197_ _23197_/A vssd1 vssd1 vccd1 vccd1 _27135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22148_ _22148_/A vssd1 vssd1 vccd1 vccd1 _22148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22079_ _22067_/X _22068_/X _22069_/X _22070_/X _22071_/X _22072_/X vssd1 vssd1 vccd1
+ vccd1 _22080_/A sky130_fd_sc_hd__mux4_1
X_26956_ _22658_/X _26956_/D vssd1 vssd1 vccd1 vccd1 _26956_/Q sky130_fd_sc_hd__dfxtp_1
X_14970_ _15708_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14970_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_965 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13921_ _13921_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _13921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25907_ _27585_/CLK _25907_/D vssd1 vssd1 vccd1 vccd1 _25907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26887_ _22412_/X _26887_/D vssd1 vssd1 vccd1 vccd1 _26887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16640_ _16640_/A vssd1 vssd1 vccd1 vccd1 _16641_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25838_ _26037_/CLK _25838_/D vssd1 vssd1 vccd1 vccd1 _25838_/Q sky130_fd_sc_hd__dfxtp_1
X_13852_ _15695_/A _15695_/C _15695_/B vssd1 vssd1 vccd1 vccd1 _14149_/B sky130_fd_sc_hd__or3b_2
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16571_ _16652_/B _16888_/B _16651_/A vssd1 vssd1 vccd1 vccd1 _16571_/X sky130_fd_sc_hd__and3b_1
X_27983__449 vssd1 vssd1 vccd1 vccd1 _27983__449/HI _27983_/A sky130_fd_sc_hd__conb_1
X_25769_ _25769_/A vssd1 vssd1 vccd1 vccd1 _27840_/D sky130_fd_sc_hd__clkbuf_1
X_13783_ _13876_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13783_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18310_ _18310_/A vssd1 vssd1 vccd1 vccd1 _25962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15522_ _15522_/A vssd1 vssd1 vccd1 vccd1 _26215_/D sky130_fd_sc_hd__clkbuf_1
X_27508_ _27511_/CLK _27508_/D vssd1 vssd1 vccd1 vccd1 _27508_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19290_ _19290_/A vssd1 vssd1 vccd1 vccd1 _19290_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _18241_/A vssd1 vssd1 vccd1 vccd1 _25959_/D sky130_fd_sc_hd__clkbuf_1
X_27439_ _27790_/CLK _27439_/D vssd1 vssd1 vccd1 vccd1 _27439_/Q sky130_fd_sc_hd__dfxtp_1
X_15453_ _15464_/A vssd1 vssd1 vccd1 vccd1 _15462_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14404_ _26654_/Q _14392_/X _14398_/X _14403_/Y vssd1 vssd1 vccd1 vccd1 _26654_/D
+ sky130_fd_sc_hd__a31o_1
X_18172_ _27806_/Q _26567_/Q _26439_/Q _26119_/Q _18099_/X _18126_/X vssd1 vssd1 vccd1
+ vccd1 _18172_/X sky130_fd_sc_hd__mux4_2
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ _14779_/X _26276_/Q _15390_/S vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17123_ _17116_/X _17117_/X _17119_/X _17122_/X vssd1 vssd1 vccd1 vccd1 _17123_/X
+ sky130_fd_sc_hd__o22a_1
X_14335_ _14335_/A _14335_/B vssd1 vssd1 vccd1 vccd1 _14335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17054_ _25916_/Q _25982_/Q _17071_/S vssd1 vssd1 vccd1 vccd1 _17055_/B sky130_fd_sc_hd__mux2_1
X_14266_ _14354_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14266_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16005_ _27481_/Q _27479_/Q _16020_/C _16004_/Y _27369_/Q vssd1 vssd1 vccd1 vccd1
+ _16112_/B sky130_fd_sc_hd__o311a_1
XFILLER_171_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13217_ _27038_/Q _13216_/X _13229_/S vssd1 vssd1 vccd1 vccd1 _13218_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14197_ _14374_/A _14200_/B vssd1 vssd1 vccd1 vccd1 _14197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _27286_/Q _13176_/B vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__and2_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _17956_/A _17813_/X vssd1 vssd1 vccd1 vccd1 _17956_/X sky130_fd_sc_hd__or2b_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _27061_/Q _13078_/X _13079_/S vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__mux2_1
Xrepeater304 _27666_/CLK vssd1 vssd1 vccd1 vccd1 _27663_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater315 _27699_/CLK vssd1 vssd1 vccd1 vccd1 _27703_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater326 _27778_/CLK vssd1 vssd1 vccd1 vccd1 _27636_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16907_ _16877_/X _16904_/Y _16906_/X vssd1 vssd1 vccd1 vccd1 _24263_/A sky130_fd_sc_hd__o21a_1
Xrepeater337 _27783_/CLK vssd1 vssd1 vccd1 vccd1 _27782_/CLK sky130_fd_sc_hd__clkbuf_1
X_17887_ _18474_/A vssd1 vssd1 vccd1 vccd1 _18479_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater348 _27669_/CLK vssd1 vssd1 vccd1 vccd1 _27667_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater359 _27585_/CLK vssd1 vssd1 vccd1 vccd1 _27348_/CLK sky130_fd_sc_hd__clkbuf_1
X_19626_ _19626_/A vssd1 vssd1 vccd1 vccd1 _19626_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16838_ _16838_/A _16838_/B vssd1 vssd1 vccd1 vccd1 _16838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19557_ _18929_/X _19556_/X _18932_/X vssd1 vssd1 vccd1 vccd1 _19557_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16769_ _16779_/A _16769_/B vssd1 vssd1 vccd1 vccd1 _16780_/A sky130_fd_sc_hd__xnor2_1
XFILLER_202_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18508_ _18502_/X _18504_/X _18507_/X _18443_/X _18489_/X vssd1 vssd1 vccd1 vccd1
+ _18509_/C sky130_fd_sc_hd__a221o_1
XFILLER_22_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19488_ _19488_/A vssd1 vssd1 vccd1 vccd1 _19488_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18439_ _18437_/X _18438_/X _18326_/X vssd1 vssd1 vccd1 vccd1 _18439_/X sky130_fd_sc_hd__o21a_1
XFILLER_194_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21450_ _21450_/A vssd1 vssd1 vccd1 vccd1 _21450_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20401_ _20401_/A vssd1 vssd1 vccd1 vccd1 _20401_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21381_ _21373_/X _21374_/X _21375_/X _21376_/X _21377_/X _21378_/X vssd1 vssd1 vccd1
+ vccd1 _21382_/A sky130_fd_sc_hd__mux4_1
XFILLER_179_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20332_ _20318_/X _20319_/X _20320_/X _20321_/X _20322_/X _20323_/X vssd1 vssd1 vccd1
+ vccd1 _20333_/A sky130_fd_sc_hd__mux4_1
X_23120_ _23120_/A vssd1 vssd1 vccd1 vccd1 _27101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23051_ _27071_/Q _17692_/X _23059_/S vssd1 vssd1 vccd1 vccd1 _23052_/A sky130_fd_sc_hd__mux2_1
X_20263_ _20263_/A vssd1 vssd1 vccd1 vccd1 _20263_/X sky130_fd_sc_hd__clkbuf_1
X_22002_ _22071_/A vssd1 vssd1 vccd1 vccd1 _22002_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20194_ _20181_/X _20183_/X _20185_/X _20187_/X _20188_/X _20189_/X vssd1 vssd1 vccd1
+ vccd1 _20195_/A sky130_fd_sc_hd__mux4_1
X_26810_ _22148_/X _26810_/D vssd1 vssd1 vccd1 vccd1 _26810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27790_ _27790_/CLK _27790_/D vssd1 vssd1 vccd1 vccd1 _27980_/A sky130_fd_sc_hd__dfxtp_1
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26741_ _21904_/X _26741_/D vssd1 vssd1 vccd1 vccd1 _26741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23953_ _23949_/X _23951_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23953_/X sky130_fd_sc_hd__mux2_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22904_ _22904_/A vssd1 vssd1 vccd1 vccd1 _22904_/X sky130_fd_sc_hd__clkbuf_1
X_26672_ _21660_/X _26672_/D vssd1 vssd1 vccd1 vccd1 _26672_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23884_ _23881_/X _23883_/X _23891_/S vssd1 vssd1 vccd1 vccd1 _23884_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25623_ _23643_/X _27981_/A _25623_/S vssd1 vssd1 vccd1 vccd1 _25624_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22835_ _22821_/X _22822_/X _22823_/X _22824_/X _22825_/X _22826_/X vssd1 vssd1 vccd1
+ vccd1 _22836_/A sky130_fd_sc_hd__mux4_1
XFILLER_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25554_ _25584_/A vssd1 vssd1 vccd1 vccd1 _25554_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22766_ _22766_/A vssd1 vssd1 vccd1 vccd1 _22766_/X sky130_fd_sc_hd__clkbuf_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24505_ _27589_/Q _24505_/B vssd1 vssd1 vccd1 vccd1 _24505_/X sky130_fd_sc_hd__or2_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ _21705_/X _21706_/X _21707_/X _21708_/X _21709_/X _21710_/X vssd1 vssd1 vccd1
+ vccd1 _21718_/A sky130_fd_sc_hd__mux4_1
XFILLER_13_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25485_ _24754_/A _25474_/X _25481_/Y _25484_/X _25467_/X vssd1 vssd1 vccd1 vccd1
+ _27761_/D sky130_fd_sc_hd__a221oi_1
XFILLER_13_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22697_ _22697_/A vssd1 vssd1 vccd1 vccd1 _22697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27224_ _27224_/CLK _27224_/D vssd1 vssd1 vccd1 vccd1 _27224_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24436_ _24480_/A vssd1 vssd1 vccd1 vccd1 _24445_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21648_ _21648_/A vssd1 vssd1 vccd1 vccd1 _21648_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27155_ _27155_/CLK _27155_/D vssd1 vssd1 vccd1 vccd1 _27155_/Q sky130_fd_sc_hd__dfxtp_1
X_24367_ _24367_/A vssd1 vssd1 vccd1 vccd1 _27465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21579_ _21579_/A vssd1 vssd1 vccd1 vccd1 _21647_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_80 _18791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_91 _19037_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26106_ _19687_/X _26106_/D vssd1 vssd1 vccd1 vccd1 _26106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_501 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23318_ _23277_/Y input57/X _27749_/Q _23301_/Y vssd1 vssd1 vccd1 vccd1 _23318_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_181_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27086_ _27294_/CLK _27086_/D vssd1 vssd1 vccd1 vccd1 _27086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24298_ _24298_/A vssd1 vssd1 vccd1 vccd1 _25618_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26037_ _26037_/CLK _26037_/D vssd1 vssd1 vccd1 vccd1 _26037_/Q sky130_fd_sc_hd__dfxtp_1
X_14051_ _26781_/Q _14042_/X _14038_/X _14050_/Y vssd1 vssd1 vccd1 vccd1 _26781_/D
+ sky130_fd_sc_hd__a31o_1
X_23249_ _23249_/A vssd1 vssd1 vccd1 vccd1 _27159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _13002_/A vssd1 vssd1 vccd1 vccd1 _27798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17810_ _18182_/A vssd1 vssd1 vccd1 vccd1 _17810_/X sky130_fd_sc_hd__clkbuf_4
X_18790_ _19412_/A vssd1 vssd1 vccd1 vccd1 _18790_/X sky130_fd_sc_hd__buf_2
XFILLER_122_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27988_ _27988_/A _15895_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17741_ _17757_/A vssd1 vssd1 vccd1 vccd1 _17754_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_48_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26939_ _22592_/X _26939_/D vssd1 vssd1 vccd1 vccd1 _26939_/Q sky130_fd_sc_hd__dfxtp_1
X_14953_ _14807_/X _26459_/Q _14955_/S vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13904_ _13904_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17672_ _17672_/A vssd1 vssd1 vccd1 vccd1 _25906_/D sky130_fd_sc_hd__clkbuf_1
X_14884_ _14884_/A vssd1 vssd1 vccd1 vccd1 _26490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19411_ _19273_/X _19410_/X _19387_/X vssd1 vssd1 vccd1 vccd1 _19411_/X sky130_fd_sc_hd__o21a_1
X_16623_ _16623_/A _16623_/B _16623_/C vssd1 vssd1 vccd1 vccd1 _16804_/A sky130_fd_sc_hd__and3_1
X_13835_ _26848_/Q _13832_/X _13833_/X _13834_/Y vssd1 vssd1 vccd1 vccd1 _26848_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_90_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19342_ _19273_/X _19341_/X _19229_/X vssd1 vssd1 vccd1 vccd1 _19342_/X sky130_fd_sc_hd__o21a_1
X_16554_ _16542_/X _16546_/X _16548_/Y _16549_/X _16553_/X vssd1 vssd1 vccd1 vccd1
+ _16554_/X sky130_fd_sc_hd__a221o_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _13857_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15505_ _15505_/A vssd1 vssd1 vccd1 vccd1 _26223_/D sky130_fd_sc_hd__clkbuf_1
X_19273_ _19431_/A vssd1 vssd1 vccd1 vccd1 _19273_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16485_ _16698_/A vssd1 vssd1 vccd1 vccd1 _16697_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13697_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13697_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ _18224_/A _17910_/X vssd1 vssd1 vccd1 vccd1 _18224_/X sky130_fd_sc_hd__or2b_1
X_15436_ _26253_/Q _13360_/X _15440_/S vssd1 vssd1 vccd1 vccd1 _15437_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18155_ _26694_/Q _26662_/Q _26630_/Q _26598_/Q _18036_/X _18106_/X vssd1 vssd1 vccd1
+ vccd1 _18157_/A sky130_fd_sc_hd__mux4_1
XFILLER_200_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15367_ _15367_/A vssd1 vssd1 vccd1 vccd1 _26284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17106_ _25920_/Q _25986_/Q _17132_/S vssd1 vssd1 vccd1 vccd1 _17107_/B sky130_fd_sc_hd__mux2_1
XFILLER_190_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14318_ _14406_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14318_/Y sky130_fd_sc_hd__nor2_1
X_18086_ _26819_/Q _26787_/Q _26755_/Q _26723_/Q _18085_/X _24388_/A vssd1 vssd1 vccd1
+ vccd1 _18086_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15298_ _26314_/Q _13369_/X _15306_/S vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17037_ _17035_/X _17036_/X _17048_/S vssd1 vssd1 vccd1 vccd1 _17037_/X sky130_fd_sc_hd__mux2_1
X_14249_ _26711_/Q _14238_/X _14242_/X _14248_/Y vssd1 vssd1 vccd1 vccd1 _26711_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _18979_/X _18981_/X _18986_/X _18866_/X _18987_/X vssd1 vssd1 vccd1 vccd1
+ _18989_/C sky130_fd_sc_hd__a221o_1
Xrepeater101 _27672_/CLK vssd1 vssd1 vccd1 vccd1 _27787_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater112 _27786_/CLK vssd1 vssd1 vccd1 vccd1 _27122_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_112_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater123 _27125_/CLK vssd1 vssd1 vccd1 vccd1 _27854_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _27596_/Q vssd1 vssd1 vccd1 vccd1 _18483_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater134 _25995_/CLK vssd1 vssd1 vccd1 vccd1 _27845_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater145 _27160_/CLK vssd1 vssd1 vccd1 vccd1 _27856_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater156 _27412_/CLK vssd1 vssd1 vccd1 vccd1 _27278_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater167 _26024_/CLK vssd1 vssd1 vccd1 vccd1 _27144_/CLK sky130_fd_sc_hd__clkbuf_1
X_20950_ _20950_/A vssd1 vssd1 vccd1 vccd1 _20950_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater178 _27109_/CLK vssd1 vssd1 vccd1 vccd1 _27110_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater189 _26013_/CLK vssd1 vssd1 vccd1 vccd1 _26014_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_26_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19609_ _19625_/A vssd1 vssd1 vccd1 vccd1 _19609_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20881_ _20864_/X _20865_/X _20866_/X _20867_/X _20870_/X _20874_/X vssd1 vssd1 vccd1
+ vccd1 _20882_/A sky130_fd_sc_hd__mux4_1
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22620_ _22620_/A vssd1 vssd1 vccd1 vccd1 _22620_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22551_ _22539_/X _22542_/X _22545_/X _22548_/X _22549_/X _22550_/X vssd1 vssd1 vccd1
+ vccd1 _22552_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21502_ _21550_/A vssd1 vssd1 vccd1 vccd1 _21502_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25270_ _25323_/A _27507_/Q vssd1 vssd1 vccd1 vccd1 _25272_/C sky130_fd_sc_hd__xnor2_1
X_22482_ _22482_/A vssd1 vssd1 vccd1 vccd1 _22482_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24221_ _25617_/A _24222_/B vssd1 vssd1 vccd1 vccd1 _27380_/D sky130_fd_sc_hd__nor2_1
X_21433_ _21427_/X _21428_/X _21429_/X _21430_/X _21431_/X _21432_/X vssd1 vssd1 vccd1
+ vccd1 _21434_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21364_ _21364_/A vssd1 vssd1 vccd1 vccd1 _21364_/X sky130_fd_sc_hd__clkbuf_1
X_24152_ _24152_/A vssd1 vssd1 vccd1 vccd1 _27348_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23103_ _27095_/Q _17769_/X _23103_/S vssd1 vssd1 vccd1 vccd1 _23104_/A sky130_fd_sc_hd__mux2_1
X_20315_ _20315_/A vssd1 vssd1 vccd1 vccd1 _20315_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21295_ _21285_/X _21286_/X _21287_/X _21288_/X _21289_/X _21290_/X vssd1 vssd1 vccd1
+ vccd1 _21296_/A sky130_fd_sc_hd__mux4_1
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24083_ _24083_/A vssd1 vssd1 vccd1 vccd1 _27317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20246_ _20232_/X _20233_/X _20234_/X _20235_/X _20236_/X _20237_/X vssd1 vssd1 vccd1
+ vccd1 _20247_/A sky130_fd_sc_hd__mux4_1
X_23034_ _23034_/A vssd1 vssd1 vccd1 vccd1 _23035_/D sky130_fd_sc_hd__inv_2
XFILLER_192_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27842_ _27842_/CLK _27842_/D vssd1 vssd1 vccd1 vccd1 _27842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20177_ _20177_/A vssd1 vssd1 vccd1 vccd1 _20177_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27773_ _27773_/CLK _27773_/D vssd1 vssd1 vccd1 vccd1 _27773_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24985_ _24982_/X _24984_/X _25003_/S vssd1 vssd1 vccd1 vccd1 _24985_/X sky130_fd_sc_hd__mux2_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26724_ _21842_/X _26724_/D vssd1 vssd1 vccd1 vccd1 _26724_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23936_ _27845_/Q _27149_/Q _25894_/Q _25862_/Q _23920_/X _23897_/X vssd1 vssd1 vccd1
+ vccd1 _23936_/X sky130_fd_sc_hd__mux4_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26655_ _21606_/X _26655_/D vssd1 vssd1 vccd1 vccd1 _26655_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23867_ _25923_/Q _25989_/Q _25822_/Q _26021_/Q _23852_/X _23835_/X vssd1 vssd1 vccd1
+ vccd1 _23867_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13620_ _26926_/Q _13613_/X _13616_/X _13619_/Y vssd1 vssd1 vccd1 vccd1 _26926_/D
+ sky130_fd_sc_hd__a31o_1
X_25606_ _24811_/A _18606_/X _25604_/X _25605_/Y _25592_/X vssd1 vssd1 vccd1 vccd1
+ _27782_/D sky130_fd_sc_hd__a221oi_1
XFILLER_199_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22818_ _22818_/A vssd1 vssd1 vccd1 vccd1 _22818_/X sky130_fd_sc_hd__clkbuf_1
X_26586_ _21366_/X _26586_/D vssd1 vssd1 vccd1 vccd1 _26586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23798_ _27070_/Q _23761_/X _23763_/X _27102_/Q _23765_/X vssd1 vssd1 vccd1 vccd1
+ _23798_/X sky130_fd_sc_hd__a221o_1
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _13923_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13551_/Y sky130_fd_sc_hd__nor2_1
X_25537_ _25530_/X _25245_/B _25536_/X _25513_/X vssd1 vssd1 vccd1 vccd1 _25537_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22749_ _22735_/X _22736_/X _22737_/X _22738_/X _22739_/X _22740_/X vssd1 vssd1 vccd1
+ vccd1 _22750_/A sky130_fd_sc_hd__mux4_1
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16270_ _16490_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16270_/Y sky130_fd_sc_hd__nor2_1
X_13482_ _13553_/A vssd1 vssd1 vccd1 vccd1 _13482_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25468_ _24744_/A _25431_/X _25460_/Y _25465_/X _25467_/X vssd1 vssd1 vccd1 vccd1
+ _27758_/D sky130_fd_sc_hd__a221oi_1
XFILLER_125_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15221_ _14753_/X _26348_/Q _15223_/S vssd1 vssd1 vccd1 vccd1 _15222_/A sky130_fd_sc_hd__mux2_1
X_27207_ _27207_/CLK _27207_/D vssd1 vssd1 vccd1 vccd1 _27207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24419_ _24419_/A vssd1 vssd1 vccd1 vccd1 _27488_/D sky130_fd_sc_hd__clkbuf_1
X_25399_ _25399_/A vssd1 vssd1 vccd1 vccd1 _27738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27138_ _27835_/CLK _27138_/D vssd1 vssd1 vccd1 vccd1 _27138_/Q sky130_fd_sc_hd__dfxtp_1
X_15152_ _15152_/A vssd1 vssd1 vccd1 vccd1 _26379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _14172_/A vssd1 vssd1 vccd1 vccd1 _14157_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15083_ _15083_/A vssd1 vssd1 vccd1 vccd1 _26410_/D sky130_fd_sc_hd__clkbuf_1
X_19960_ _19976_/A vssd1 vssd1 vccd1 vccd1 _19960_/X sky130_fd_sc_hd__clkbuf_2
X_27069_ _27415_/CLK _27069_/D vssd1 vssd1 vccd1 vccd1 _27069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14034_ _26786_/Q _14024_/X _14019_/X _14033_/Y vssd1 vssd1 vccd1 vccd1 _26786_/D
+ sky130_fd_sc_hd__a31o_1
X_18911_ _19501_/A _18911_/B vssd1 vssd1 vccd1 vccd1 _18911_/X sky130_fd_sc_hd__or2_1
XFILLER_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19891_ _19891_/A vssd1 vssd1 vccd1 vccd1 _19891_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18842_ _18842_/A _18842_/B _18842_/C vssd1 vssd1 vccd1 vccd1 _18843_/A sky130_fd_sc_hd__and3_1
XFILLER_121_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18773_ _18945_/A vssd1 vssd1 vccd1 vccd1 _19296_/S sky130_fd_sc_hd__clkbuf_2
X_15985_ _15985_/A vssd1 vssd1 vccd1 vccd1 _15985_/Y sky130_fd_sc_hd__inv_2
X_27989__455 vssd1 vssd1 vccd1 vccd1 _27989__455/HI _27989_/A sky130_fd_sc_hd__conb_1
X_17724_ _27423_/Q vssd1 vssd1 vccd1 vccd1 _17724_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14936_ _14782_/X _26467_/Q _14940_/S vssd1 vssd1 vccd1 vccd1 _14937_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17655_ _17655_/A vssd1 vssd1 vccd1 vccd1 _25898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ _14867_/A vssd1 vssd1 vccd1 vccd1 _26498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13818_ _26854_/Q _13806_/X _13807_/X _13817_/Y vssd1 vssd1 vccd1 vccd1 _26854_/D
+ sky130_fd_sc_hd__a31o_1
X_16606_ _16392_/Y _16399_/Y _16433_/Y vssd1 vssd1 vccd1 vccd1 _16606_/Y sky130_fd_sc_hd__o21ai_1
X_17586_ _17586_/A vssd1 vssd1 vccd1 vccd1 _17595_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14798_ _14798_/A vssd1 vssd1 vccd1 vccd1 _14798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19325_ _19316_/X _19319_/X _19323_/X _19324_/X _19258_/X vssd1 vssd1 vccd1 vccd1
+ _19336_/B sky130_fd_sc_hd__a221o_1
X_16537_ _27396_/Q _16312_/X _16412_/X _25964_/Q _16536_/Y vssd1 vssd1 vccd1 vccd1
+ _16822_/A sky130_fd_sc_hd__a221o_2
X_13749_ _26879_/Q _13737_/X _13745_/X _13748_/Y vssd1 vssd1 vccd1 vccd1 _26879_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19256_ _27810_/Q _26571_/Q _26443_/Q _26123_/Q _19255_/X _19183_/X vssd1 vssd1 vccd1
+ vccd1 _19256_/X sky130_fd_sc_hd__mux4_2
X_16468_ _16768_/B vssd1 vssd1 vccd1 vccd1 _16611_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18207_ _18322_/A vssd1 vssd1 vccd1 vccd1 _18207_/X sky130_fd_sc_hd__clkbuf_1
X_15419_ _15419_/A vssd1 vssd1 vccd1 vccd1 _26261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19187_ _19178_/X _19181_/X _19185_/X _19186_/X _19139_/X vssd1 vssd1 vccd1 vccd1
+ _19201_/B sky130_fd_sc_hd__a221o_1
X_16399_ _16383_/A _16393_/Y _16397_/X _16398_/X vssd1 vssd1 vccd1 vccd1 _16399_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_191_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18138_ _18138_/A _18066_/X vssd1 vssd1 vccd1 vccd1 _18138_/X sky130_fd_sc_hd__or2b_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18069_ _26274_/Q _26242_/Q _26210_/Q _26178_/Q _18044_/X _18068_/X vssd1 vssd1 vccd1
+ vccd1 _18069_/X sky130_fd_sc_hd__mux4_2
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20100_ _20272_/A vssd1 vssd1 vccd1 vccd1 _20165_/A sky130_fd_sc_hd__buf_2
XFILLER_99_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21080_ _21128_/A vssd1 vssd1 vccd1 vccd1 _21080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20031_ _20079_/A vssd1 vssd1 vccd1 vccd1 _20031_/X sky130_fd_sc_hd__clkbuf_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24770_ _27622_/Q _24758_/X _24769_/Y _24760_/X vssd1 vssd1 vccd1 vccd1 _27622_/D
+ sky130_fd_sc_hd__o211a_1
X_21982_ _21998_/A vssd1 vssd1 vccd1 vccd1 _21982_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23721_ _23721_/A vssd1 vssd1 vccd1 vccd1 _27264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20933_ _20921_/X _20922_/X _20923_/X _20924_/X _20925_/X _20926_/X vssd1 vssd1 vccd1
+ vccd1 _20934_/A sky130_fd_sc_hd__mux4_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26440_ _20855_/X _26440_/D vssd1 vssd1 vccd1 vccd1 _26440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23652_ _23720_/S vssd1 vssd1 vccd1 vccd1 _23661_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20864_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20864_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22603_ _22593_/X _22594_/X _22595_/X _22596_/X _22597_/X _22598_/X vssd1 vssd1 vccd1
+ vccd1 _22604_/A sky130_fd_sc_hd__mux4_1
X_26371_ _20609_/X _26371_/D vssd1 vssd1 vccd1 vccd1 _26371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23583_ _23583_/A vssd1 vssd1 vccd1 vccd1 _27215_/D sky130_fd_sc_hd__clkbuf_1
X_20795_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20795_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25322_ _27715_/Q _25308_/X _25321_/Y _25297_/X vssd1 vssd1 vccd1 vccd1 _27715_/D
+ sky130_fd_sc_hd__o211a_1
X_22534_ _22534_/A vssd1 vssd1 vccd1 vccd1 _22534_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25253_ _25261_/A _25253_/B vssd1 vssd1 vccd1 vccd1 _25253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22465_ _22452_/X _22454_/X _22456_/X _22458_/X _22459_/X _22460_/X vssd1 vssd1 vccd1
+ vccd1 _22466_/A sky130_fd_sc_hd__mux4_1
XFILLER_183_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24204_ _24298_/A vssd1 vssd1 vccd1 vccd1 _24217_/A sky130_fd_sc_hd__buf_4
XFILLER_120_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21416_ _21464_/A vssd1 vssd1 vccd1 vccd1 _21416_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25184_ _25308_/A vssd1 vssd1 vccd1 vccd1 _25184_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22396_ _22396_/A vssd1 vssd1 vccd1 vccd1 _22396_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24135_ _24135_/A vssd1 vssd1 vccd1 vccd1 _27340_/D sky130_fd_sc_hd__clkbuf_1
X_21347_ _21341_/X _21342_/X _21343_/X _21344_/X _21345_/X _21346_/X vssd1 vssd1 vccd1
+ vccd1 _21348_/A sky130_fd_sc_hd__mux4_1
XFILLER_120_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24066_ _27383_/Q _24072_/B vssd1 vssd1 vccd1 vccd1 _24067_/A sky130_fd_sc_hd__and2_1
X_21278_ _21278_/A vssd1 vssd1 vccd1 vccd1 _21278_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23017_ _23009_/X _23010_/X _23011_/X _23012_/X _23013_/X _23014_/X vssd1 vssd1 vccd1
+ vccd1 _23018_/A sky130_fd_sc_hd__mux4_1
XFILLER_150_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20229_ _20229_/A vssd1 vssd1 vccd1 vccd1 _20229_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27825_ _27825_/CLK _27825_/D vssd1 vssd1 vccd1 vccd1 _27825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15770_ _26111_/Q _15760_/X _15766_/X _15769_/Y vssd1 vssd1 vccd1 vccd1 _26111_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12982_/A vssd1 vssd1 vccd1 vccd1 _27807_/D sky130_fd_sc_hd__clkbuf_1
X_27756_ _27756_/CLK _27756_/D vssd1 vssd1 vccd1 vccd1 _27756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24968_ _27670_/Q _24838_/A _24967_/Y _24663_/A vssd1 vssd1 vccd1 vccd1 _27670_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14721_ _14721_/A vssd1 vssd1 vccd1 vccd1 _14721_/X sky130_fd_sc_hd__buf_2
X_26707_ _21788_/X _26707_/D vssd1 vssd1 vccd1 vccd1 _26707_/Q sky130_fd_sc_hd__dfxtp_1
X_23919_ _23896_/X _23917_/X _23918_/X _23911_/X vssd1 vssd1 vccd1 vccd1 _27287_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27687_ _27791_/CLK _27687_/D vssd1 vssd1 vccd1 vccd1 _27978_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24899_ _24913_/A _24899_/B vssd1 vssd1 vccd1 vccd1 _24899_/Y sky130_fd_sc_hd__nand2_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ _27413_/Q vssd1 vssd1 vccd1 vccd1 _17440_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26638_ _21542_/X _26638_/D vssd1 vssd1 vccd1 vccd1 _26638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _26576_/Q _14645_/X _14640_/X _14651_/Y vssd1 vssd1 vccd1 vccd1 _26576_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13603_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ _17338_/X _17371_/B vssd1 vssd1 vccd1 vccd1 _17371_/X sky130_fd_sc_hd__and2b_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _26601_/Q _14576_/X _14579_/X _14582_/Y vssd1 vssd1 vccd1 vccd1 _26601_/D
+ sky130_fd_sc_hd__a31o_1
X_26569_ _21300_/X _26569_/D vssd1 vssd1 vccd1 vccd1 _26569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19110_ _19460_/A vssd1 vssd1 vccd1 vccd1 _19407_/A sky130_fd_sc_hd__buf_4
XFILLER_14_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16322_ _16353_/A vssd1 vssd1 vccd1 vccd1 _16490_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_201_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13534_ _26949_/Q _13510_/X _13528_/X _13533_/Y vssd1 vssd1 vccd1 vccd1 _26949_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1012 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19041_ _19113_/A _19041_/B vssd1 vssd1 vccd1 vccd1 _19041_/X sky130_fd_sc_hd__or2_1
X_16253_ _27391_/Q _16132_/A _16137_/X _26057_/Q _16252_/X vssd1 vssd1 vccd1 vccd1
+ _24290_/A sky130_fd_sc_hd__a221o_1
X_13465_ _27360_/Q _13062_/A _13082_/A _27328_/Q _13092_/X vssd1 vssd1 vccd1 vccd1
+ _16298_/A sky130_fd_sc_hd__a221oi_4
X_15204_ _14727_/X _26356_/Q _15212_/S vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16184_ _27376_/Q _16244_/B _16244_/C vssd1 vssd1 vccd1 vccd1 _16184_/X sky130_fd_sc_hd__and3_1
XFILLER_138_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _26978_/Q _13395_/X _13399_/S vssd1 vssd1 vccd1 vccd1 _13397_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15135_ _15135_/A vssd1 vssd1 vccd1 vccd1 _26387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19943_ _19991_/A vssd1 vssd1 vccd1 vccd1 _19943_/X sky130_fd_sc_hd__clkbuf_1
X_15066_ _14737_/X _26417_/Q _15068_/S vssd1 vssd1 vccd1 vccd1 _15067_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14017_ _14383_/A _14029_/B vssd1 vssd1 vccd1 vccd1 _14017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19874_ _19866_/X _19867_/X _19868_/X _19869_/X _19870_/X _19871_/X vssd1 vssd1 vccd1
+ vccd1 _19875_/A sky130_fd_sc_hd__mux4_1
X_18825_ _18897_/A vssd1 vssd1 vccd1 vccd1 _19399_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18756_ _18756_/A vssd1 vssd1 vccd1 vccd1 _26038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15968_ _15980_/A vssd1 vssd1 vccd1 vccd1 _15973_/A sky130_fd_sc_hd__buf_2
XFILLER_83_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17707_ _17707_/A vssd1 vssd1 vccd1 vccd1 _25921_/D sky130_fd_sc_hd__clkbuf_1
X_14919_ _14919_/A vssd1 vssd1 vccd1 vccd1 _26475_/D sky130_fd_sc_hd__clkbuf_1
X_15899_ _15899_/A vssd1 vssd1 vccd1 vccd1 _15899_/Y sky130_fd_sc_hd__inv_2
X_18687_ _26008_/Q _17772_/X _18689_/S vssd1 vssd1 vccd1 vccd1 _18688_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ _17638_/A vssd1 vssd1 vccd1 vccd1 _25890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ _17479_/X _25860_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17570_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19308_ _26541_/Q _26509_/Q _26477_/Q _27053_/Q _19297_/X _19407_/A vssd1 vssd1 vccd1
+ vccd1 _19308_/X sky130_fd_sc_hd__mux4_1
X_20580_ _20566_/X _20567_/X _20568_/X _20569_/X _20570_/X _20571_/X vssd1 vssd1 vccd1
+ vccd1 _20581_/A sky130_fd_sc_hd__mux4_1
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19239_ _19191_/X _19238_/X _19194_/X vssd1 vssd1 vccd1 vccd1 _19239_/X sky130_fd_sc_hd__o21a_1
XFILLER_143_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22250_ _22250_/A vssd1 vssd1 vccd1 vccd1 _22250_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21201_ _21195_/X _21196_/X _21197_/X _21198_/X _21199_/X _21200_/X vssd1 vssd1 vccd1
+ vccd1 _21202_/A sky130_fd_sc_hd__mux4_1
X_22181_ _22525_/A vssd1 vssd1 vccd1 vccd1 _22250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21132_ _21200_/A vssd1 vssd1 vccd1 vccd1 _21132_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25940_ _27149_/CLK _25940_/D vssd1 vssd1 vccd1 vccd1 _25940_/Q sky130_fd_sc_hd__dfxtp_1
X_21063_ _21149_/A vssd1 vssd1 vccd1 vccd1 _21128_/A sky130_fd_sc_hd__buf_2
XFILLER_115_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20014_ _20272_/A vssd1 vssd1 vccd1 vccd1 _20079_/A sky130_fd_sc_hd__buf_2
X_25871_ _27157_/CLK _25871_/D vssd1 vssd1 vccd1 vccd1 _25871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24822_ _27639_/Q _24813_/X _24821_/Y _24817_/X vssd1 vssd1 vccd1 vccd1 _27639_/D
+ sky130_fd_sc_hd__o211a_1
X_27610_ _27610_/CLK _27610_/D vssd1 vssd1 vccd1 vccd1 _27610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27541_ _27541_/CLK _27541_/D vssd1 vssd1 vccd1 vccd1 _27541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24753_ _27615_/Q _24742_/X _24752_/Y _24746_/X vssd1 vssd1 vccd1 vccd1 _27615_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _21997_/A vssd1 vssd1 vccd1 vccd1 _21965_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23704_ _23704_/A vssd1 vssd1 vccd1 vccd1 _27256_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20916_/A vssd1 vssd1 vccd1 vccd1 _20916_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27472_ _27472_/CLK _27472_/D vssd1 vssd1 vccd1 vccd1 _27472_/Q sky130_fd_sc_hd__dfxtp_1
X_24684_ _16979_/B _24673_/X _24683_/X _24677_/X vssd1 vssd1 vccd1 vccd1 _27591_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21896_ _21912_/A vssd1 vssd1 vccd1 vccd1 _21896_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_508 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26423_ _20785_/X _26423_/D vssd1 vssd1 vccd1 vccd1 _26423_/Q sky130_fd_sc_hd__dfxtp_1
X_23635_ _23638_/A _23638_/C _23634_/Y vssd1 vssd1 vccd1 vccd1 _27229_/D sky130_fd_sc_hd__o21a_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _20847_/A vssd1 vssd1 vccd1 vccd1 _20847_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26354_ _20549_/X _26354_/D vssd1 vssd1 vccd1 vccd1 _26354_/Q sky130_fd_sc_hd__dfxtp_1
X_23566_ _23566_/A vssd1 vssd1 vccd1 vccd1 _27210_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20778_ _20770_/X _20771_/X _20772_/X _20773_/X _20775_/X _20777_/X vssd1 vssd1 vccd1
+ vccd1 _20779_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25305_ _25329_/A _25329_/B vssd1 vssd1 vccd1 vccd1 _25306_/B sky130_fd_sc_hd__xnor2_2
X_22517_ _22503_/X _22504_/X _22505_/X _22506_/X _22507_/X _22508_/X vssd1 vssd1 vccd1
+ vccd1 _22518_/A sky130_fd_sc_hd__mux4_1
XFILLER_168_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26285_ _20309_/X _26285_/D vssd1 vssd1 vccd1 vccd1 _26285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23497_ _27192_/Q _23500_/B vssd1 vssd1 vccd1 vccd1 _23497_/X sky130_fd_sc_hd__or2_1
XFILLER_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25236_ _25266_/B _25242_/B vssd1 vssd1 vccd1 vccd1 _25237_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ _27033_/Q _13038_/X _13258_/S vssd1 vssd1 vccd1 vccd1 _13251_/A sky130_fd_sc_hd__mux2_1
X_22448_ _22448_/A vssd1 vssd1 vccd1 vccd1 _22448_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25167_ _27696_/Q _25142_/X _25166_/Y _25132_/X vssd1 vssd1 vccd1 vccd1 _27696_/D
+ sky130_fd_sc_hd__o211a_1
X_13181_ _13181_/A vssd1 vssd1 vccd1 vccd1 _27044_/D sky130_fd_sc_hd__clkbuf_1
X_22379_ _22366_/X _22368_/X _22370_/X _22372_/X _22373_/X _22374_/X vssd1 vssd1 vccd1
+ vccd1 _22380_/A sky130_fd_sc_hd__mux4_1
XFILLER_159_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24118_ _24118_/A vssd1 vssd1 vccd1 vccd1 _27333_/D sky130_fd_sc_hd__clkbuf_1
X_25098_ _25098_/A vssd1 vssd1 vccd1 vccd1 _27686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24049_ _23849_/A _24047_/X _24048_/X _23864_/A vssd1 vssd1 vccd1 vccd1 _27302_/D
+ sky130_fd_sc_hd__o211a_1
X_16940_ _27601_/Q vssd1 vssd1 vccd1 vccd1 _19448_/A sky130_fd_sc_hd__inv_2
XFILLER_111_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16871_ _27575_/Q _24218_/A _25615_/A vssd1 vssd1 vccd1 vccd1 _16872_/D sky130_fd_sc_hd__and3_1
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18610_ _27541_/Q _27520_/Q vssd1 vssd1 vccd1 vccd1 _18610_/X sky130_fd_sc_hd__and2_1
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27808_ _25682_/X _27808_/D vssd1 vssd1 vccd1 vccd1 _27808_/Q sky130_fd_sc_hd__dfxtp_1
X_15822_ _15822_/A vssd1 vssd1 vccd1 vccd1 _26089_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19590_ _19638_/A vssd1 vssd1 vccd1 vccd1 _19590_/X sky130_fd_sc_hd__clkbuf_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15753_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18541_ _18437_/X _18540_/X _18483_/X vssd1 vssd1 vccd1 vccd1 _18541_/X sky130_fd_sc_hd__o21a_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _27814_/Q _12965_/B vssd1 vssd1 vccd1 vccd1 _12966_/A sky130_fd_sc_hd__and2_1
X_27739_ _27750_/CLK _27739_/D vssd1 vssd1 vccd1 vccd1 _27739_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _26556_/Q _14698_/X _14693_/X _14703_/Y vssd1 vssd1 vccd1 vccd1 _26556_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18472_ _26836_/Q _26804_/Q _26772_/Q _26740_/Q _18358_/X _18380_/X vssd1 vssd1 vccd1
+ vccd1 _18472_/X sky130_fd_sc_hd__mux4_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ _15684_/A vssd1 vssd1 vccd1 vccd1 _26143_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 _13331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _15708_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14635_/Y sky130_fd_sc_hd__nor2_1
X_17423_ _24061_/A _17674_/B _17601_/C vssd1 vssd1 vccd1 vccd1 _17505_/A sky130_fd_sc_hd__or3_2
XANTENNA_362 _27407_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_373 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 _25641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _17299_/X _17349_/X _17351_/X _17353_/X vssd1 vssd1 vccd1 vccd1 _17354_/X
+ sky130_fd_sc_hd__o22a_1
X_14566_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14566_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13517_ _13904_/A _13517_/B vssd1 vssd1 vccd1 vccd1 _13517_/Y sky130_fd_sc_hd__nor2_1
X_16305_ _16125_/B _16304_/B _16639_/A vssd1 vssd1 vccd1 vccd1 _16603_/A sky130_fd_sc_hd__a21o_1
XFILLER_202_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17285_ _17283_/X _17284_/X _17296_/S vssd1 vssd1 vccd1 vccd1 _17285_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ _14497_/A vssd1 vssd1 vccd1 vccd1 _15756_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19024_ _19014_/X _19017_/X _19021_/X _19022_/X _19023_/X vssd1 vssd1 vccd1 vccd1
+ _19037_/B sky130_fd_sc_hd__a221o_2
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16236_ _27528_/Q _15992_/A vssd1 vssd1 vccd1 vccd1 _16236_/X sky130_fd_sc_hd__or2b_1
XFILLER_173_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13448_ _13868_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16167_ _27386_/Q vssd1 vssd1 vccd1 vccd1 _16426_/A sky130_fd_sc_hd__inv_2
X_13379_ _14769_/A vssd1 vssd1 vccd1 vccd1 _13379_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _15407_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15175_/A sky130_fd_sc_hd__nor2_4
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16098_ _16098_/A vssd1 vssd1 vccd1 vccd1 _16098_/X sky130_fd_sc_hd__buf_2
XFILLER_170_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19926_ _20272_/A vssd1 vssd1 vccd1 vccd1 _19991_/A sky130_fd_sc_hd__clkbuf_2
X_15049_ _14709_/X _26425_/Q _15057_/S vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19857_ _19857_/A vssd1 vssd1 vccd1 vccd1 _19857_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18808_ _18828_/A vssd1 vssd1 vccd1 vccd1 _19401_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19788_ _19780_/X _19781_/X _19782_/X _19783_/X _19784_/X _19785_/X vssd1 vssd1 vccd1
+ vccd1 _19789_/A sky130_fd_sc_hd__mux4_1
XFILLER_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18739_ _18739_/A vssd1 vssd1 vccd1 vccd1 _26030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21750_ _21750_/A vssd1 vssd1 vccd1 vccd1 _21750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20701_ _20701_/A vssd1 vssd1 vccd1 vccd1 _20701_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21681_ _21667_/X _21670_/X _21673_/X _21676_/X _21677_/X _21678_/X vssd1 vssd1 vccd1
+ vccd1 _21682_/A sky130_fd_sc_hd__mux4_1
XFILLER_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23420_ _23598_/A vssd1 vssd1 vccd1 vccd1 _23624_/A sky130_fd_sc_hd__buf_2
X_20632_ _20617_/X _20619_/X _20621_/X _20623_/X _20624_/X _20625_/X vssd1 vssd1 vccd1
+ vccd1 _20633_/A sky130_fd_sc_hd__mux4_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23351_ _24844_/A _27238_/Q vssd1 vssd1 vccd1 vccd1 _23351_/Y sky130_fd_sc_hd__xnor2_1
X_20563_ _20563_/A vssd1 vssd1 vccd1 vccd1 _20563_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22302_ _22350_/A vssd1 vssd1 vccd1 vccd1 _22302_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26070_ _26073_/CLK _26070_/D vssd1 vssd1 vccd1 vccd1 _26070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23282_ _27731_/Q input42/X vssd1 vssd1 vccd1 vccd1 _23282_/X sky130_fd_sc_hd__xor2_1
XFILLER_34_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20494_ _20480_/X _20481_/X _20482_/X _20483_/X _20484_/X _20485_/X vssd1 vssd1 vccd1
+ vccd1 _20495_/A sky130_fd_sc_hd__mux4_1
XFILLER_118_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25021_ _25019_/X _25020_/X _25046_/S vssd1 vssd1 vccd1 vccd1 _25021_/X sky130_fd_sc_hd__mux2_1
X_22233_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22164_ _22164_/A vssd1 vssd1 vccd1 vccd1 _22164_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21115_ _21109_/X _21110_/X _21111_/X _21112_/X _21113_/X _21114_/X vssd1 vssd1 vccd1
+ vccd1 _21116_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22095_ _22083_/X _22084_/X _22085_/X _22086_/X _22088_/X _22090_/X vssd1 vssd1 vccd1
+ vccd1 _22096_/A sky130_fd_sc_hd__mux4_1
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26972_ _22710_/X _26972_/D vssd1 vssd1 vccd1 vccd1 _26972_/Q sky130_fd_sc_hd__dfxtp_1
X_25923_ _25923_/CLK _25923_/D vssd1 vssd1 vccd1 vccd1 _25923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21046_ _21114_/A vssd1 vssd1 vccd1 vccd1 _21046_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_530 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25854_ _25989_/CLK _25854_/D vssd1 vssd1 vccd1 vccd1 _25854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24805_ _27634_/Q _24798_/X _24804_/Y _24801_/X vssd1 vssd1 vccd1 vccd1 _27634_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25785_ _25785_/A vssd1 vssd1 vccd1 vccd1 _27847_/D sky130_fd_sc_hd__clkbuf_1
X_22997_ _23029_/A vssd1 vssd1 vccd1 vccd1 _22997_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27524_ _27529_/CLK _27524_/D vssd1 vssd1 vccd1 vccd1 _27524_/Q sky130_fd_sc_hd__dfxtp_1
X_24736_ _24803_/A vssd1 vssd1 vccd1 vccd1 _24970_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_21948_ _21948_/A vssd1 vssd1 vccd1 vccd1 _21948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_828 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27455_ _27458_/CLK _27455_/D vssd1 vssd1 vccd1 vccd1 _27455_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24667_ _27169_/Q _24671_/B vssd1 vssd1 vccd1 vccd1 _24667_/X sky130_fd_sc_hd__or2_1
X_21879_ _21911_/A vssd1 vssd1 vccd1 vccd1 _21879_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14420_ _26649_/Q _14405_/X _14416_/X _14419_/Y vssd1 vssd1 vccd1 vccd1 _26649_/D
+ sky130_fd_sc_hd__a31o_1
X_26406_ _20731_/X _26406_/D vssd1 vssd1 vccd1 vccd1 _26406_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23618_ _23618_/A vssd1 vssd1 vccd1 vccd1 _27224_/D sky130_fd_sc_hd__clkbuf_1
X_27386_ _27386_/CLK _27386_/D vssd1 vssd1 vccd1 vccd1 _27386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24598_ _27659_/Q _24598_/B vssd1 vssd1 vccd1 vccd1 _24599_/A sky130_fd_sc_hd__and2_1
XFILLER_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14351_ _26674_/Q _14337_/X _14345_/X _14350_/Y vssd1 vssd1 vccd1 vccd1 _26674_/D
+ sky130_fd_sc_hd__a31o_1
X_26337_ _20491_/X _26337_/D vssd1 vssd1 vccd1 vccd1 _26337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23549_ _23549_/A vssd1 vssd1 vccd1 vccd1 _27205_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _27009_/Q _13198_/X _13302_/S vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__mux2_1
X_17070_ _27831_/Q _27135_/Q _25880_/Q _25848_/Q _17015_/X _17069_/X vssd1 vssd1 vccd1
+ vccd1 _17070_/X sky130_fd_sc_hd__mux4_1
X_14282_ _26699_/Q _14270_/X _14271_/X _14281_/Y vssd1 vssd1 vccd1 vccd1 _26699_/D
+ sky130_fd_sc_hd__a31o_1
X_26268_ _20245_/X _26268_/D vssd1 vssd1 vccd1 vccd1 _26268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16021_ _16030_/A _16030_/B _16030_/C _16020_/X vssd1 vssd1 vccd1 vccd1 _16205_/A
+ sky130_fd_sc_hd__nor4b_1
X_28007_ _28007_/A _15859_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_25219_ _25212_/A _25211_/B _25211_/A vssd1 vssd1 vccd1 vccd1 _25220_/B sky130_fd_sc_hd__a21boi_1
X_13233_ _16177_/A vssd1 vssd1 vccd1 vccd1 _14807_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26199_ _20007_/X _26199_/D vssd1 vssd1 vccd1 vccd1 _26199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13164_ _27283_/Q _13201_/B vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__and2_2
XFILLER_123_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17972_ _18150_/A vssd1 vssd1 vccd1 vccd1 _17972_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13095_ _27059_/Q _13094_/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13096_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19711_ _19727_/A vssd1 vssd1 vccd1 vccd1 _19711_/X sky130_fd_sc_hd__clkbuf_1
X_16923_ _25572_/A _25582_/A _25583_/A _25584_/A _25108_/A vssd1 vssd1 vccd1 vccd1
+ _18584_/A sky130_fd_sc_hd__o311a_1
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19642_ _22613_/A vssd1 vssd1 vccd1 vccd1 _25725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16854_ _16625_/A _16764_/A _16395_/A _16625_/B vssd1 vssd1 vccd1 vccd1 _16854_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _13111_/X _26096_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15806_/A sky130_fd_sc_hd__mux2_1
X_19573_ _19834_/A vssd1 vssd1 vccd1 vccd1 _19639_/A sky130_fd_sc_hd__clkbuf_2
X_13997_ _26796_/Q _13987_/X _13983_/X _13996_/Y vssd1 vssd1 vccd1 vccd1 _26796_/D
+ sky130_fd_sc_hd__a31o_1
X_16785_ _16785_/A _16785_/B vssd1 vssd1 vccd1 vccd1 _16785_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18524_ _18524_/A _17799_/X vssd1 vssd1 vccd1 vccd1 _18524_/X sky130_fd_sc_hd__or2b_1
X_15736_ _15736_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15736_/Y sky130_fd_sc_hd__nor2_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ _27821_/Q _12952_/B vssd1 vssd1 vccd1 vccd1 _12949_/A sky130_fd_sc_hd__and2_1
XFILLER_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18455_ _18455_/A vssd1 vssd1 vccd1 vccd1 _18455_/X sky130_fd_sc_hd__buf_2
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_170 _16033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15667_ _13166_/X _26150_/Q _15667_/S vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__mux2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _14464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_192 _16451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17406_ _17406_/A vssd1 vssd1 vccd1 vccd1 _17407_/A sky130_fd_sc_hd__buf_2
X_14618_ _15779_/A _14620_/B vssd1 vssd1 vccd1 vccd1 _14618_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18386_ _18311_/X _18378_/X _18385_/X _18253_/X vssd1 vssd1 vccd1 vccd1 _18398_/B
+ sky130_fd_sc_hd__a211o_1
X_15598_ _26181_/Q _14775_/A _15606_/S vssd1 vssd1 vccd1 vccd1 _15599_/A sky130_fd_sc_hd__mux2_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17337_ _27853_/Q _27157_/Q _25902_/Q _25870_/Q _17325_/X _17313_/X vssd1 vssd1 vccd1
+ vccd1 _17337_/X sky130_fd_sc_hd__mux4_1
X_14549_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14549_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17268_ _17216_/X _17268_/B vssd1 vssd1 vccd1 vccd1 _17268_/X sky130_fd_sc_hd__and2b_1
XFILLER_88_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19007_ _26400_/Q _26368_/Q _26336_/Q _26304_/Q _18887_/X _18982_/X vssd1 vssd1 vccd1
+ vccd1 _19007_/X sky130_fd_sc_hd__mux4_1
X_16219_ _27523_/Q _15991_/A vssd1 vssd1 vccd1 vccd1 _16219_/X sky130_fd_sc_hd__or2b_1
X_17199_ _17197_/X _17198_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19909_ _19909_/A vssd1 vssd1 vccd1 vccd1 _19909_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22920_ _22920_/A vssd1 vssd1 vccd1 vccd1 _22920_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22851_ _22837_/X _22838_/X _22839_/X _22840_/X _22841_/X _22842_/X vssd1 vssd1 vccd1
+ vccd1 _22852_/A sky130_fd_sc_hd__mux4_1
XFILLER_72_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21802_ _21802_/A vssd1 vssd1 vccd1 vccd1 _21802_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25570_ _27711_/Q _25568_/X _25569_/X vssd1 vssd1 vccd1 vccd1 _25570_/Y sky130_fd_sc_hd__a21oi_1
X_22782_ _22782_/A vssd1 vssd1 vccd1 vccd1 _22782_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24521_ _24551_/S vssd1 vssd1 vccd1 vccd1 _24631_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_21733_ _21721_/X _21722_/X _21723_/X _21724_/X _21725_/X _21726_/X vssd1 vssd1 vccd1
+ vccd1 _21734_/A sky130_fd_sc_hd__mux4_1
XFILLER_197_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27240_ _27245_/CLK _27240_/D vssd1 vssd1 vccd1 vccd1 _27240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24452_ _27624_/Q _24456_/B vssd1 vssd1 vccd1 vccd1 _24453_/A sky130_fd_sc_hd__and2_1
XFILLER_61_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21664_ _21664_/A vssd1 vssd1 vccd1 vccd1 _21664_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23403_ _24756_/A _27242_/Q _27252_/Q _24782_/A _23402_/X vssd1 vssd1 vccd1 vccd1
+ _23409_/C sky130_fd_sc_hd__a221o_1
X_20615_ _20615_/A vssd1 vssd1 vccd1 vccd1 _20615_/X sky130_fd_sc_hd__clkbuf_1
X_27171_ _27587_/CLK _27171_/D vssd1 vssd1 vccd1 vccd1 _27171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24383_ _25524_/A vssd1 vssd1 vccd1 vccd1 _24384_/A sky130_fd_sc_hd__clkbuf_2
X_21595_ _21580_/X _21582_/X _21584_/X _21586_/X _21587_/X _21588_/X vssd1 vssd1 vccd1
+ vccd1 _21596_/A sky130_fd_sc_hd__mux4_1
X_26122_ _19739_/X _26122_/D vssd1 vssd1 vccd1 vccd1 _26122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23334_ _27237_/Q vssd1 vssd1 vccd1 vccd1 _23334_/Y sky130_fd_sc_hd__inv_2
X_20546_ _20531_/X _20533_/X _20535_/X _20537_/X _20538_/X _20539_/X vssd1 vssd1 vccd1
+ vccd1 _20547_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26053_ _26053_/CLK _26053_/D vssd1 vssd1 vccd1 vccd1 _26053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23265_ _23260_/Y input71/X _27748_/Q _23261_/Y _23264_/X vssd1 vssd1 vccd1 vccd1
+ _23275_/B sky130_fd_sc_hd__a221o_1
XFILLER_134_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20477_ _20477_/A vssd1 vssd1 vccd1 vccd1 _20477_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25004_ _27069_/Q _27101_/Q _25004_/S vssd1 vssd1 vccd1 vccd1 _25004_/X sky130_fd_sc_hd__mux2_1
X_22216_ _22264_/A vssd1 vssd1 vccd1 vccd1 _22216_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23196_ _17440_/X _27135_/Q _23204_/S vssd1 vssd1 vccd1 vccd1 _23197_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22147_ _22141_/X _22142_/X _22143_/X _22144_/X _22145_/X _22146_/X vssd1 vssd1 vccd1
+ vccd1 _22148_/A sky130_fd_sc_hd__mux4_1
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_688 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22078_ _22078_/A vssd1 vssd1 vccd1 vccd1 _22078_/X sky130_fd_sc_hd__clkbuf_1
X_26955_ _22656_/X _26955_/D vssd1 vssd1 vccd1 vccd1 _26955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13920_ _13920_/A vssd1 vssd1 vccd1 vccd1 _13930_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25906_ _27857_/CLK _25906_/D vssd1 vssd1 vccd1 vccd1 _25906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21029_ _21023_/X _21024_/X _21025_/X _21026_/X _21027_/X _21028_/X vssd1 vssd1 vccd1
+ vccd1 _21030_/A sky130_fd_sc_hd__mux4_1
X_26886_ _22410_/X _26886_/D vssd1 vssd1 vccd1 vccd1 _26886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13851_ _16017_/B vssd1 vssd1 vccd1 vccd1 _15695_/B sky130_fd_sc_hd__clkbuf_1
X_25837_ _27851_/CLK _25837_/D vssd1 vssd1 vccd1 vccd1 _25837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13782_ _26868_/Q _13778_/X _13780_/X _13781_/Y vssd1 vssd1 vccd1 vccd1 _26868_/D
+ sky130_fd_sc_hd__a31o_1
X_16570_ _16648_/C _16570_/B vssd1 vssd1 vccd1 vccd1 _16651_/A sky130_fd_sc_hd__nand2_1
X_25768_ _17469_/X _27840_/Q _25768_/S vssd1 vssd1 vccd1 vccd1 _25769_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15521_ _13161_/X _26215_/Q _15523_/S vssd1 vssd1 vccd1 vccd1 _15522_/A sky130_fd_sc_hd__mux2_1
X_27507_ _27629_/CLK _27507_/D vssd1 vssd1 vccd1 vccd1 _27507_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24719_ _27188_/Q _24725_/B vssd1 vssd1 vccd1 vccd1 _24719_/X sky130_fd_sc_hd__or2_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25699_ _25689_/X _25690_/X _25691_/X _25692_/X _25693_/X _25694_/X vssd1 vssd1 vccd1
+ vccd1 _25700_/A sky130_fd_sc_hd__mux4_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15452_ _15452_/A vssd1 vssd1 vccd1 vccd1 _26246_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18240_ _18264_/A _18240_/B _18240_/C vssd1 vssd1 vccd1 vccd1 _18241_/A sky130_fd_sc_hd__and3_1
X_27438_ _27672_/CLK _27438_/D vssd1 vssd1 vccd1 vccd1 _27438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_494 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14403_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14403_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15383_ _15383_/A vssd1 vssd1 vccd1 vccd1 _26277_/D sky130_fd_sc_hd__clkbuf_1
X_18171_ _18171_/A vssd1 vssd1 vccd1 vccd1 _25956_/D sky130_fd_sc_hd__clkbuf_1
X_27369_ _27576_/CLK _27369_/D vssd1 vssd1 vccd1 vccd1 _27369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14334_ _26680_/Q _14322_/X _14329_/X _14333_/Y vssd1 vssd1 vccd1 vccd1 _26680_/D
+ sky130_fd_sc_hd__a31o_1
X_17122_ _17120_/X _17121_/X _17098_/X vssd1 vssd1 vccd1 vccd1 _17122_/X sky130_fd_sc_hd__a21bo_1
XFILLER_51_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17053_ _27830_/Q _27134_/Q _25879_/Q _25847_/Q _17015_/X _16989_/X vssd1 vssd1 vccd1
+ vccd1 _17053_/X sky130_fd_sc_hd__mux4_1
X_14265_ _14304_/A vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16004_ _27483_/Q _27374_/Q vssd1 vssd1 vccd1 vccd1 _16004_/Y sky130_fd_sc_hd__xnor2_1
X_13216_ _14798_/A vssd1 vssd1 vccd1 vccd1 _13216_/X sky130_fd_sc_hd__buf_2
XFILLER_87_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14196_ _26730_/Q _14186_/X _14194_/X _14195_/Y vssd1 vssd1 vccd1 vccd1 _26730_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13147_/A vssd1 vssd1 vccd1 vccd1 _27050_/D sky130_fd_sc_hd__clkbuf_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17955_ _26686_/Q _26654_/Q _26622_/Q _26590_/Q _17865_/X _17928_/X vssd1 vssd1 vccd1
+ vccd1 _17956_/A sky130_fd_sc_hd__mux4_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13078_ _14724_/A vssd1 vssd1 vccd1 vccd1 _13078_/X sky130_fd_sc_hd__buf_2
Xrepeater305 _27668_/CLK vssd1 vssd1 vccd1 vccd1 _27666_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater316 _27695_/CLK vssd1 vssd1 vccd1 vccd1 _27699_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16836_/A _16598_/A _16647_/X _16905_/X vssd1 vssd1 vccd1 vccd1 _16906_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater327 _27250_/CLK vssd1 vssd1 vccd1 vccd1 _27778_/CLK sky130_fd_sc_hd__clkbuf_1
X_17886_ _17884_/X _17885_/X _17886_/S vssd1 vssd1 vccd1 vccd1 _17886_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater338 _27784_/CLK vssd1 vssd1 vccd1 vccd1 _27783_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater349 _27645_/CLK vssd1 vssd1 vccd1 vccd1 _27669_/CLK sky130_fd_sc_hd__clkbuf_1
X_19625_ _19625_/A vssd1 vssd1 vccd1 vccd1 _19625_/X sky130_fd_sc_hd__clkbuf_2
X_16837_ _16835_/Y _16599_/A _16793_/D _16598_/A _16836_/Y vssd1 vssd1 vccd1 vccd1
+ _16838_/B sky130_fd_sc_hd__a32o_1
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19556_ _26841_/Q _26809_/Q _26777_/Q _26745_/Q _18778_/X _18930_/X vssd1 vssd1 vccd1
+ vccd1 _19556_/X sky130_fd_sc_hd__mux4_2
XFILLER_202_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ _16783_/A _16768_/B vssd1 vssd1 vccd1 vccd1 _16768_/X sky130_fd_sc_hd__xor2_1
XFILLER_202_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18507_ _18505_/X _18506_/X _18580_/S vssd1 vssd1 vccd1 vccd1 _18507_/X sky130_fd_sc_hd__mux2_2
X_15719_ _26130_/Q _15705_/X _15713_/X _15718_/Y vssd1 vssd1 vccd1 vccd1 _26130_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19487_ _26293_/Q _26261_/Q _26229_/Q _26197_/Q _19441_/X _19486_/X vssd1 vssd1 vccd1
+ vccd1 _19487_/X sky130_fd_sc_hd__mux4_1
X_16699_ _16699_/A _16808_/B vssd1 vssd1 vccd1 vccd1 _16699_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18438_ _26290_/Q _26258_/Q _26226_/Q _26194_/Q _18301_/X _18324_/X vssd1 vssd1 vccd1
+ vccd1 _18438_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18369_ _18369_/A _17799_/X vssd1 vssd1 vccd1 vccd1 _18369_/X sky130_fd_sc_hd__or2b_1
XFILLER_147_522 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20400_ _20392_/X _20393_/X _20394_/X _20395_/X _20396_/X _20397_/X vssd1 vssd1 vccd1
+ vccd1 _20401_/A sky130_fd_sc_hd__mux4_1
X_21380_ _21380_/A vssd1 vssd1 vccd1 vccd1 _21380_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20331_ _20331_/A vssd1 vssd1 vccd1 vccd1 _20331_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23050_ _23107_/S vssd1 vssd1 vccd1 vccd1 _23059_/S sky130_fd_sc_hd__clkbuf_2
X_20262_ _20248_/X _20249_/X _20250_/X _20251_/X _20253_/X _20255_/X vssd1 vssd1 vccd1
+ vccd1 _20263_/A sky130_fd_sc_hd__mux4_1
X_22001_ _22087_/A vssd1 vssd1 vccd1 vccd1 _22071_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20193_ _20193_/A vssd1 vssd1 vccd1 vccd1 _20193_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26740_ _21902_/X _26740_/D vssd1 vssd1 vccd1 vccd1 _26740_/Q sky130_fd_sc_hd__dfxtp_1
X_23952_ _27788_/Q vssd1 vssd1 vccd1 vccd1 _23987_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22903_ _22888_/X _22890_/X _22892_/X _22894_/X _22895_/X _22896_/X vssd1 vssd1 vccd1
+ vccd1 _22904_/A sky130_fd_sc_hd__mux4_1
X_26671_ _21658_/X _26671_/D vssd1 vssd1 vccd1 vccd1 _26671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_553 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23883_ _25925_/Q _25991_/Q _25824_/Q _26023_/Q _23852_/X _23882_/X vssd1 vssd1 vccd1
+ vccd1 _23883_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25622_ _25622_/A vssd1 vssd1 vccd1 vccd1 _27790_/D sky130_fd_sc_hd__clkbuf_1
X_22834_ _22834_/A vssd1 vssd1 vccd1 vccd1 _22834_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25553_ _25553_/A vssd1 vssd1 vccd1 vccd1 _25553_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_197_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22765_ _22751_/X _22752_/X _22753_/X _22754_/X _22755_/X _22756_/X vssd1 vssd1 vccd1
+ vccd1 _22766_/A sky130_fd_sc_hd__mux4_1
XFILLER_169_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24504_ _24405_/A _24633_/C _24503_/X _24499_/X vssd1 vssd1 vccd1 vccd1 _27522_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21716_ _21716_/A vssd1 vssd1 vccd1 vccd1 _21716_/X sky130_fd_sc_hd__clkbuf_1
X_25484_ _25470_/X _25174_/B _25482_/X _25483_/X vssd1 vssd1 vccd1 vccd1 _25484_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22696_ _22696_/A vssd1 vssd1 vccd1 vccd1 _22696_/X sky130_fd_sc_hd__clkbuf_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24435_ _24435_/A vssd1 vssd1 vccd1 vccd1 _24480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27223_ _27224_/CLK _27223_/D vssd1 vssd1 vccd1 vccd1 _27223_/Q sky130_fd_sc_hd__dfxtp_1
X_21647_ _21647_/A vssd1 vssd1 vccd1 vccd1 _21647_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27154_ _27154_/CLK _27154_/D vssd1 vssd1 vccd1 vccd1 _27154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24366_ _27565_/Q _24372_/B vssd1 vssd1 vccd1 vccd1 _24367_/A sky130_fd_sc_hd__and2_1
XFILLER_197_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21578_ _21578_/A vssd1 vssd1 vccd1 vccd1 _21578_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_70 _18402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 _18796_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26105_ _19685_/X _26105_/D vssd1 vssd1 vccd1 vccd1 _26105_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_92 _19046_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23317_ _27728_/Q _23315_/Y _23312_/Y input54/X _23316_/X vssd1 vssd1 vccd1 vccd1
+ _23320_/C sky130_fd_sc_hd__a221o_1
X_27085_ _27786_/CLK _27085_/D vssd1 vssd1 vccd1 vccd1 _27085_/Q sky130_fd_sc_hd__dfxtp_1
X_20529_ _20529_/A vssd1 vssd1 vccd1 vccd1 _20529_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24297_ _24297_/A _24302_/B vssd1 vssd1 vccd1 vccd1 _27428_/D sky130_fd_sc_hd__nor2_1
XFILLER_119_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26036_ _27851_/CLK _26036_/D vssd1 vssd1 vccd1 vccd1 _26036_/Q sky130_fd_sc_hd__dfxtp_1
X_14050_ _14406_/A _14060_/B vssd1 vssd1 vccd1 vccd1 _14050_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23248_ _17517_/X _27159_/Q _23248_/S vssd1 vssd1 vccd1 vccd1 _23249_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13001_ _27798_/Q _13009_/B vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__and2_1
XFILLER_134_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23179_ _23179_/A vssd1 vssd1 vccd1 vccd1 _27128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27987_ _27987_/A _15896_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
XFILLER_47_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17740_ _27428_/Q vssd1 vssd1 vccd1 vccd1 _17740_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26938_ _22590_/X _26938_/D vssd1 vssd1 vccd1 vccd1 _26938_/Q sky130_fd_sc_hd__dfxtp_1
X_14952_ _14952_/A vssd1 vssd1 vccd1 vccd1 _26460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13903_ _26825_/Q _13893_/X _13899_/X _13902_/Y vssd1 vssd1 vccd1 vccd1 _26825_/D
+ sky130_fd_sc_hd__a31o_1
X_17671_ _17523_/X _25906_/Q _17671_/S vssd1 vssd1 vccd1 vccd1 _17672_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26869_ _22346_/X _26869_/D vssd1 vssd1 vccd1 vccd1 _26869_/Q sky130_fd_sc_hd__dfxtp_1
X_14883_ _26490_/Q _13420_/X _14883_/S vssd1 vssd1 vccd1 vccd1 _14884_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19410_ _26706_/Q _26674_/Q _26642_/Q _26610_/Q _19317_/X _19385_/X vssd1 vssd1 vccd1
+ vccd1 _19410_/X sky130_fd_sc_hd__mux4_1
X_16622_ _16559_/A _16623_/B _16535_/A vssd1 vssd1 vccd1 vccd1 _16804_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13834_ _13926_/A _13838_/B vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19341_ _26703_/Q _26671_/Q _26639_/Q _26607_/Q _19317_/X _19227_/X vssd1 vssd1 vccd1
+ vccd1 _19341_/X sky130_fd_sc_hd__mux4_2
X_13765_ _13779_/A vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16553_ _16550_/X _16551_/Y _16552_/Y vssd1 vssd1 vccd1 vccd1 _16553_/X sky130_fd_sc_hd__o21a_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15504_ _13116_/X _26223_/Q _15512_/S vssd1 vssd1 vccd1 vccd1 _15505_/A sky130_fd_sc_hd__mux2_1
X_19272_ _19409_/A _19272_/B vssd1 vssd1 vccd1 vccd1 _19272_/X sky130_fd_sc_hd__or2_1
XFILLER_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13696_ _26899_/Q _13682_/X _13692_/X _13695_/Y vssd1 vssd1 vccd1 vccd1 _26899_/D
+ sky130_fd_sc_hd__a31o_1
X_16484_ _16446_/Y _16447_/Y _16460_/Y _16255_/Y _25910_/Q vssd1 vssd1 vccd1 vccd1
+ _16497_/B sky130_fd_sc_hd__a41o_1
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18223_ _26697_/Q _26665_/Q _26633_/Q _26601_/Q _18004_/X _18005_/X vssd1 vssd1 vccd1
+ vccd1 _18224_/A sky130_fd_sc_hd__mux4_2
X_15435_ _15435_/A vssd1 vssd1 vccd1 vccd1 _26254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18154_ _26822_/Q _26790_/Q _26758_/Q _26726_/Q _18034_/X _18058_/X vssd1 vssd1 vccd1
+ vccd1 _18154_/X sky130_fd_sc_hd__mux4_1
X_15366_ _14753_/X _26284_/Q _15368_/S vssd1 vssd1 vccd1 vccd1 _15367_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17105_ _27834_/Q _27138_/Q _25883_/Q _25851_/Q _17081_/X _17069_/X vssd1 vssd1 vccd1
+ vccd1 _17105_/X sky130_fd_sc_hd__mux4_1
X_14317_ _26686_/Q _14310_/X _14311_/X _14316_/Y vssd1 vssd1 vccd1 vccd1 _26686_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18085_ _18085_/A vssd1 vssd1 vccd1 vccd1 _18085_/X sky130_fd_sc_hd__clkbuf_4
X_15297_ _15319_/A vssd1 vssd1 vccd1 vccd1 _15306_/S sky130_fd_sc_hd__clkbuf_2
X_14248_ _14335_/A _14248_/B vssd1 vssd1 vccd1 vccd1 _14248_/Y sky130_fd_sc_hd__nor2_1
X_17036_ _27068_/Q _27100_/Q _17047_/S vssd1 vssd1 vccd1 vccd1 _17036_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _14356_/A _14187_/B vssd1 vssd1 vccd1 vccd1 _14179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _19220_/A vssd1 vssd1 vccd1 vccd1 _18987_/X sky130_fd_sc_hd__clkbuf_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater102 _25901_/CLK vssd1 vssd1 vccd1 vccd1 _27852_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater113 _27288_/CLK vssd1 vssd1 vccd1 vccd1 _27786_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _26269_/Q _26237_/Q _26205_/Q _26173_/Q _17873_/X _17937_/X vssd1 vssd1 vccd1
+ vccd1 _17938_/X sky130_fd_sc_hd__mux4_1
XFILLER_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater124 _26037_/CLK vssd1 vssd1 vccd1 vccd1 _27855_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater135 _25996_/CLK vssd1 vssd1 vccd1 vccd1 _25995_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater146 _27160_/CLK vssd1 vssd1 vccd1 vccd1 _27211_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater157 _27412_/CLK vssd1 vssd1 vccd1 vccd1 _27408_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater168 _27081_/CLK vssd1 vssd1 vccd1 vccd1 _26024_/CLK sky130_fd_sc_hd__clkbuf_1
X_17869_ _17779_/X _17862_/X _17868_/X _24396_/A vssd1 vssd1 vccd1 vccd1 _17881_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater179 _27096_/CLK vssd1 vssd1 vccd1 vccd1 _27109_/CLK sky130_fd_sc_hd__clkbuf_1
X_19608_ _19640_/A vssd1 vssd1 vccd1 vccd1 _19608_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20880_ _20880_/A vssd1 vssd1 vccd1 vccd1 _20880_/X sky130_fd_sc_hd__clkbuf_1
X_19539_ _19537_/X _19538_/X _19539_/S vssd1 vssd1 vccd1 vccd1 _19539_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22550_ _22598_/A vssd1 vssd1 vccd1 vccd1 _22550_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21501_ _21549_/A vssd1 vssd1 vccd1 vccd1 _21501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22481_ _22471_/X _22472_/X _22473_/X _22474_/X _22475_/X _22476_/X vssd1 vssd1 vccd1
+ vccd1 _22482_/A sky130_fd_sc_hd__mux4_1
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24220_ _25616_/A _24222_/B vssd1 vssd1 vccd1 vccd1 _27379_/D sky130_fd_sc_hd__nor2_1
X_21432_ _21464_/A vssd1 vssd1 vccd1 vccd1 _21432_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24151_ _27453_/Q _24151_/B vssd1 vssd1 vccd1 vccd1 _24152_/A sky130_fd_sc_hd__and2_1
XFILLER_163_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21363_ _21357_/X _21358_/X _21359_/X _21360_/X _21361_/X _21362_/X vssd1 vssd1 vccd1
+ vccd1 _21364_/A sky130_fd_sc_hd__mux4_1
XFILLER_147_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23102_ _23102_/A vssd1 vssd1 vccd1 vccd1 _27094_/D sky130_fd_sc_hd__clkbuf_1
X_20314_ _20302_/X _20303_/X _20304_/X _20305_/X _20306_/X _20307_/X vssd1 vssd1 vccd1
+ vccd1 _20315_/A sky130_fd_sc_hd__mux4_1
X_24082_ _27390_/Q _24084_/B vssd1 vssd1 vccd1 vccd1 _24083_/A sky130_fd_sc_hd__and2_1
X_21294_ _21294_/A vssd1 vssd1 vccd1 vccd1 _21294_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23033_ _23033_/A _27380_/Q _27377_/Q _27376_/Q vssd1 vssd1 vccd1 vccd1 _23034_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20245_ _20245_/A vssd1 vssd1 vccd1 vccd1 _20245_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27841_ _27842_/CLK _27841_/D vssd1 vssd1 vccd1 vccd1 _27841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20176_ _20162_/X _20163_/X _20164_/X _20165_/X _20167_/X _20169_/X vssd1 vssd1 vccd1
+ vccd1 _20177_/A sky130_fd_sc_hd__mux4_1
XFILLER_67_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27772_ _27772_/CLK _27772_/D vssd1 vssd1 vccd1 vccd1 _27772_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24984_ _25913_/Q _25979_/Q _25812_/Q _26011_/Q _24974_/X _24983_/X vssd1 vssd1 vccd1
+ vccd1 _24984_/X sky130_fd_sc_hd__mux4_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26723_ _21840_/X _26723_/D vssd1 vssd1 vccd1 vccd1 _26723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23935_ _23896_/X _23933_/X _23934_/X _23911_/X vssd1 vssd1 vccd1 vccd1 _27289_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26654_ _21598_/X _26654_/D vssd1 vssd1 vccd1 vccd1 _26654_/Q sky130_fd_sc_hd__dfxtp_1
X_23866_ _27837_/Q _27141_/Q _25886_/Q _25854_/Q _23826_/X _23850_/X vssd1 vssd1 vccd1
+ vccd1 _23866_/X sky130_fd_sc_hd__mux4_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25605_ _27718_/Q _25433_/X _25435_/X vssd1 vssd1 vccd1 vccd1 _25605_/Y sky130_fd_sc_hd__a21oi_1
X_22817_ _22802_/X _22804_/X _22806_/X _22808_/X _22809_/X _22810_/X vssd1 vssd1 vccd1
+ vccd1 _22818_/A sky130_fd_sc_hd__mux4_1
XFILLER_77_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26585_ _21364_/X _26585_/D vssd1 vssd1 vccd1 vccd1 _26585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23797_ _23795_/X _23796_/X _23797_/S vssd1 vssd1 vccd1 vccd1 _23797_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13550_ _14507_/A vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__buf_2
XFILLER_41_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25536_ _25517_/X _25522_/X _25523_/X _24904_/B _25524_/X vssd1 vssd1 vccd1 vccd1
+ _25536_/X sky130_fd_sc_hd__o311a_1
X_22748_ _22748_/A vssd1 vssd1 vccd1 vccd1 _22748_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13481_ _26960_/Q _13464_/X _13457_/X _13480_/Y vssd1 vssd1 vccd1 vccd1 _26960_/D
+ sky130_fd_sc_hd__a31o_1
X_25467_ _25592_/A vssd1 vssd1 vccd1 vccd1 _25467_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22679_ _22665_/X _22666_/X _22667_/X _22668_/X _22669_/X _22670_/X vssd1 vssd1 vccd1
+ vccd1 _22680_/A sky130_fd_sc_hd__mux4_1
XFILLER_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ _15220_/A vssd1 vssd1 vccd1 vccd1 _26349_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24418_ _27589_/Q _24422_/B vssd1 vssd1 vccd1 vccd1 _24419_/A sky130_fd_sc_hd__and2_1
X_27206_ _27208_/CLK _27206_/D vssd1 vssd1 vccd1 vccd1 _27206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25398_ _27738_/Q input49/X _25402_/S vssd1 vssd1 vccd1 vccd1 _25399_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15151_ _26379_/Q _13366_/X _15151_/S vssd1 vssd1 vccd1 vccd1 _15152_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24349_ _24349_/A vssd1 vssd1 vccd1 vccd1 _27457_/D sky130_fd_sc_hd__clkbuf_1
X_27137_ _27835_/CLK _27137_/D vssd1 vssd1 vccd1 vccd1 _27137_/Q sky130_fd_sc_hd__dfxtp_1
X_14102_ _26764_/Q _14090_/X _14093_/X _14101_/Y vssd1 vssd1 vccd1 vccd1 _26764_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_844 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15082_ _14759_/X _26410_/Q _15090_/S vssd1 vssd1 vccd1 vccd1 _15083_/A sky130_fd_sc_hd__mux2_1
X_27068_ _27677_/CLK _27068_/D vssd1 vssd1 vccd1 vccd1 _27068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ _14394_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14033_/Y sky130_fd_sc_hd__nor2_1
X_18910_ _26685_/Q _26653_/Q _26621_/Q _26589_/Q _18908_/X _18909_/X vssd1 vssd1 vccd1
+ vccd1 _18911_/B sky130_fd_sc_hd__mux4_1
X_26019_ _27417_/CLK _26019_/D vssd1 vssd1 vccd1 vccd1 _26019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19890_ _19882_/X _19883_/X _19884_/X _19885_/X _19886_/X _19887_/X vssd1 vssd1 vccd1
+ vccd1 _19891_/A sky130_fd_sc_hd__mux4_1
XFILLER_45_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18841_ _18812_/X _18822_/X _18835_/X _18837_/X _18840_/X vssd1 vssd1 vccd1 vccd1
+ _18842_/C sky130_fd_sc_hd__a221o_1
XFILLER_122_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_626 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18772_ _18969_/A _18772_/B vssd1 vssd1 vccd1 vccd1 _18772_/X sky130_fd_sc_hd__or2_1
XFILLER_121_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15984_ _15985_/A vssd1 vssd1 vccd1 vccd1 _15984_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17723_ _17723_/A vssd1 vssd1 vccd1 vccd1 _25926_/D sky130_fd_sc_hd__clkbuf_1
X_14935_ _14935_/A vssd1 vssd1 vccd1 vccd1 _26468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17654_ _17498_/X _25898_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _17655_/A sky130_fd_sc_hd__mux2_1
X_14866_ _26498_/Q _13395_/X _14868_/S vssd1 vssd1 vccd1 vccd1 _14867_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16605_ _16602_/A _16088_/Y _16093_/X _16604_/Y vssd1 vssd1 vccd1 vccd1 _25572_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_13817_ _13910_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17585_ _17585_/A vssd1 vssd1 vccd1 vccd1 _25867_/D sky130_fd_sc_hd__clkbuf_1
X_14797_ _14797_/A vssd1 vssd1 vccd1 vccd1 _26527_/D sky130_fd_sc_hd__clkbuf_1
X_19324_ _19324_/A vssd1 vssd1 vccd1 vccd1 _19324_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16536_ _16536_/A _16536_/B vssd1 vssd1 vccd1 vccd1 _16536_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13748_ _13928_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13748_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19255_ _19414_/A vssd1 vssd1 vccd1 vccd1 _19255_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_32_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16467_ _16779_/B _16441_/B _16466_/X vssd1 vssd1 vccd1 vccd1 _16692_/B sky130_fd_sc_hd__a21boi_1
XFILLER_188_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13679_ _26905_/Q _13665_/X _13676_/X _13678_/Y vssd1 vssd1 vccd1 vccd1 _26905_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18206_ _26152_/Q _26088_/Q _27016_/Q _26984_/Q _18182_/X _18112_/X vssd1 vssd1 vccd1
+ vccd1 _18208_/A sky130_fd_sc_hd__mux4_1
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15418_ _26261_/Q _13334_/X _15418_/S vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__mux2_1
X_19186_ _19324_/A vssd1 vssd1 vccd1 vccd1 _19186_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16398_ _16751_/B _16398_/B vssd1 vssd1 vccd1 vccd1 _16398_/X sky130_fd_sc_hd__and2_1
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18137_ _26149_/Q _26085_/Q _27013_/Q _26981_/Q _18041_/X _18112_/X vssd1 vssd1 vccd1
+ vccd1 _18138_/A sky130_fd_sc_hd__mux4_1
XFILLER_172_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15349_ _14727_/X _26292_/Q _15357_/S vssd1 vssd1 vccd1 vccd1 _15350_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18068_ _18324_/A vssd1 vssd1 vccd1 vccd1 _18068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17019_ _25913_/Q _25979_/Q _17071_/S vssd1 vssd1 vccd1 vccd1 _17020_/B sky130_fd_sc_hd__mux2_1
XFILLER_160_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20030_ _20078_/A vssd1 vssd1 vccd1 vccd1 _20030_/X sky130_fd_sc_hd__clkbuf_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_987 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21981_ _21997_/A vssd1 vssd1 vccd1 vccd1 _21981_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23720_ _27784_/Q _27264_/Q _23720_/S vssd1 vssd1 vccd1 vccd1 _23721_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20932_ _20932_/A vssd1 vssd1 vccd1 vccd1 _20932_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23651_ _23707_/A vssd1 vssd1 vccd1 vccd1 _23720_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_199_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20863_ _20863_/A vssd1 vssd1 vccd1 vccd1 _20863_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22602_ _22602_/A vssd1 vssd1 vccd1 vccd1 _22602_/X sky130_fd_sc_hd__clkbuf_1
X_26370_ _20607_/X _26370_/D vssd1 vssd1 vccd1 vccd1 _26370_/Q sky130_fd_sc_hd__dfxtp_1
X_23582_ _23596_/A _23582_/B vssd1 vssd1 vccd1 vccd1 _23583_/A sky130_fd_sc_hd__and2_1
X_20794_ _21145_/A vssd1 vssd1 vccd1 vccd1 _20865_/A sky130_fd_sc_hd__clkbuf_2
X_25321_ _25344_/A _25321_/B vssd1 vssd1 vccd1 vccd1 _25321_/Y sky130_fd_sc_hd__nand2_1
X_22533_ _22519_/X _22520_/X _22521_/X _22522_/X _22524_/X _22526_/X vssd1 vssd1 vccd1
+ vccd1 _22534_/A sky130_fd_sc_hd__mux4_1
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25252_ _25265_/A _25252_/B vssd1 vssd1 vccd1 vccd1 _25253_/B sky130_fd_sc_hd__xor2_1
X_22464_ _22464_/A vssd1 vssd1 vccd1 vccd1 _22464_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24203_ _25733_/A _25625_/S vssd1 vssd1 vccd1 vccd1 _24298_/A sky130_fd_sc_hd__or2_1
X_21415_ _21463_/A vssd1 vssd1 vccd1 vccd1 _21415_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25183_ _27698_/Q _25142_/X _25182_/Y _25175_/X vssd1 vssd1 vccd1 vccd1 _27698_/D
+ sky130_fd_sc_hd__o211a_1
X_22395_ _22385_/X _22386_/X _22387_/X _22388_/X _22389_/X _22390_/X vssd1 vssd1 vccd1
+ vccd1 _22396_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24134_ _27445_/Q _24140_/B vssd1 vssd1 vccd1 vccd1 _24135_/A sky130_fd_sc_hd__and2_1
XFILLER_68_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21346_ _21378_/A vssd1 vssd1 vccd1 vccd1 _21346_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24065_ _24065_/A vssd1 vssd1 vccd1 vccd1 _27309_/D sky130_fd_sc_hd__clkbuf_1
X_21277_ _21269_/X _21270_/X _21271_/X _21272_/X _21273_/X _21274_/X vssd1 vssd1 vccd1
+ vccd1 _21278_/A sky130_fd_sc_hd__mux4_1
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23016_ _23016_/A vssd1 vssd1 vccd1 vccd1 _23016_/X sky130_fd_sc_hd__clkbuf_1
X_20228_ _20216_/X _20217_/X _20218_/X _20219_/X _20220_/X _20221_/X vssd1 vssd1 vccd1
+ vccd1 _20229_/A sky130_fd_sc_hd__mux4_1
XFILLER_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_486 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27824_ _25732_/X _27824_/D vssd1 vssd1 vccd1 vccd1 _27824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ _20159_/A vssd1 vssd1 vccd1 vccd1 _20159_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _27807_/Q _12987_/B vssd1 vssd1 vccd1 vccd1 _12982_/A sky130_fd_sc_hd__and2_1
XFILLER_18_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27755_ _27756_/CLK _27755_/D vssd1 vssd1 vccd1 vccd1 _27755_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24967_ _24970_/A _24967_/B vssd1 vssd1 vccd1 vccd1 _24967_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26706_ _21786_/X _26706_/D vssd1 vssd1 vccd1 vccd1 _26706_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14720_ _14720_/A vssd1 vssd1 vccd1 vccd1 _26551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23918_ _27082_/Q _23907_/X _23908_/X _27114_/Q _23909_/X vssd1 vssd1 vccd1 vccd1
+ _23918_/X sky130_fd_sc_hd__a221o_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27686_ _27686_/CLK _27686_/D vssd1 vssd1 vccd1 vccd1 _27977_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24898_ _24902_/B _24898_/B vssd1 vssd1 vccd1 vccd1 _24899_/B sky130_fd_sc_hd__or2_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26637_ _21540_/X _26637_/D vssd1 vssd1 vccd1 vccd1 _26637_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14651_ _15725_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23849_ _23849_/A vssd1 vssd1 vccd1 vccd1 _23849_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13602_ _13602_/A vssd1 vssd1 vccd1 vccd1 _13656_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _25942_/Q _26008_/Q _17370_/S vssd1 vssd1 vccd1 vccd1 _17371_/B sky130_fd_sc_hd__mux2_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _15743_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14582_/Y sky130_fd_sc_hd__nor2_1
X_26568_ _21298_/X _26568_/D vssd1 vssd1 vccd1 vccd1 _26568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16321_ _16384_/A vssd1 vssd1 vccd1 vccd1 _16501_/A sky130_fd_sc_hd__clkbuf_2
X_13533_ _13913_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13533_/Y sky130_fd_sc_hd__nor2_1
X_25519_ _25500_/X _25221_/B _25518_/X _25513_/X vssd1 vssd1 vccd1 vccd1 _25519_/X
+ sky130_fd_sc_hd__a211o_1
X_26499_ _21056_/X _26499_/D vssd1 vssd1 vccd1 vccd1 _26499_/Q sky130_fd_sc_hd__dfxtp_1
X_19040_ _26818_/Q _26786_/Q _26754_/Q _26722_/Q _19039_/X _18967_/X vssd1 vssd1 vccd1
+ vccd1 _19041_/B sky130_fd_sc_hd__mux4_1
XFILLER_199_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13464_ _13558_/A vssd1 vssd1 vccd1 vccd1 _13464_/X sky130_fd_sc_hd__clkbuf_2
X_16252_ _16252_/A _16252_/B _16252_/C vssd1 vssd1 vccd1 vccd1 _16252_/X sky130_fd_sc_hd__and3_1
XFILLER_174_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ _15260_/S vssd1 vssd1 vccd1 vccd1 _15212_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _14785_/A vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_12_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16183_ _16194_/C vssd1 vssd1 vccd1 vccd1 _16221_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_5_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15134_ _26387_/Q _13341_/X _15140_/S vssd1 vssd1 vccd1 vccd1 _15135_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19942_ _19990_/A vssd1 vssd1 vccd1 vccd1 _19942_/X sky130_fd_sc_hd__clkbuf_1
X_15065_ _15065_/A vssd1 vssd1 vccd1 vccd1 _26418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14016_ _16442_/A vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19873_ _19873_/A vssd1 vssd1 vccd1 vccd1 _19873_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18824_ _19343_/A vssd1 vssd1 vccd1 vccd1 _18824_/X sky130_fd_sc_hd__buf_4
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18755_ _26038_/Q _17766_/X _18757_/S vssd1 vssd1 vccd1 vccd1 _18756_/A sky130_fd_sc_hd__mux2_1
X_15967_ _15967_/A vssd1 vssd1 vccd1 vccd1 _15967_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17706_ _25921_/Q _17705_/X _17706_/S vssd1 vssd1 vccd1 vccd1 _17707_/A sky130_fd_sc_hd__mux2_1
X_14918_ _14756_/X _26475_/Q _14918_/S vssd1 vssd1 vccd1 vccd1 _14919_/A sky130_fd_sc_hd__mux2_1
X_18686_ _18686_/A vssd1 vssd1 vccd1 vccd1 _26007_/D sky130_fd_sc_hd__clkbuf_1
X_15898_ _15899_/A vssd1 vssd1 vccd1 vccd1 _15898_/Y sky130_fd_sc_hd__inv_2
X_17637_ _17472_/X _25890_/Q _17645_/S vssd1 vssd1 vccd1 vccd1 _17638_/A sky130_fd_sc_hd__mux2_1
X_14849_ _26506_/Q _13369_/X _14857_/S vssd1 vssd1 vccd1 vccd1 _14850_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17568_ _17568_/A vssd1 vssd1 vccd1 vccd1 _25859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19307_ _26413_/Q _26381_/Q _26349_/Q _26317_/Q _19297_/X _19407_/A vssd1 vssd1 vccd1
+ vccd1 _19307_/X sky130_fd_sc_hd__mux4_1
X_16519_ _16824_/A _16519_/B vssd1 vssd1 vccd1 vccd1 _16550_/B sky130_fd_sc_hd__xnor2_1
X_17499_ _17498_/X _25834_/Q _17502_/S vssd1 vssd1 vccd1 vccd1 _17500_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19238_ _26282_/Q _26250_/Q _26218_/Q _26186_/Q _19144_/X _19192_/X vssd1 vssd1 vccd1
+ vccd1 _19238_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19169_ _19073_/X _19168_/X _19076_/X vssd1 vssd1 vccd1 vccd1 _19169_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21200_ _21200_/A vssd1 vssd1 vccd1 vccd1 _21200_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22180_ _22616_/A vssd1 vssd1 vccd1 vccd1 _22525_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21131_ _21217_/A vssd1 vssd1 vccd1 vccd1 _21200_/A sky130_fd_sc_hd__buf_2
XFILLER_132_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21062_ _21127_/A vssd1 vssd1 vccd1 vccd1 _21062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20013_ _20078_/A vssd1 vssd1 vccd1 vccd1 _20013_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25870_ _27157_/CLK _25870_/D vssd1 vssd1 vccd1 vccd1 _25870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24821_ _24969_/A _25601_/B vssd1 vssd1 vccd1 vccd1 _24821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27540_ _27541_/CLK _27540_/D vssd1 vssd1 vccd1 vccd1 _27540_/Q sky130_fd_sc_hd__dfxtp_1
X_21964_ _21964_/A vssd1 vssd1 vccd1 vccd1 _21964_/X sky130_fd_sc_hd__clkbuf_1
X_24752_ _24752_/A _24759_/B vssd1 vssd1 vccd1 vccd1 _24752_/Y sky130_fd_sc_hd__nand2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23703_ _27776_/Q _27256_/Q _23705_/S vssd1 vssd1 vccd1 vccd1 _23704_/A sky130_fd_sc_hd__mux2_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20915_ _20905_/X _20906_/X _20907_/X _20908_/X _20909_/X _20910_/X vssd1 vssd1 vccd1
+ vccd1 _20916_/A sky130_fd_sc_hd__mux4_1
XFILLER_199_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24683_ _27175_/Q _24685_/B vssd1 vssd1 vccd1 vccd1 _24683_/X sky130_fd_sc_hd__or2_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27471_ _27542_/CLK _27471_/D vssd1 vssd1 vccd1 vccd1 _27471_/Q sky130_fd_sc_hd__dfxtp_1
X_21895_ _21911_/A vssd1 vssd1 vccd1 vccd1 _21895_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23634_ _23638_/A _23638_/C _25430_/B vssd1 vssd1 vccd1 vccd1 _23634_/Y sky130_fd_sc_hd__a21oi_1
X_26422_ _20783_/X _26422_/D vssd1 vssd1 vccd1 vccd1 _26422_/Q sky130_fd_sc_hd__dfxtp_1
X_20846_ _20832_/X _20833_/X _20834_/X _20835_/X _20836_/X _20837_/X vssd1 vssd1 vccd1
+ vccd1 _20847_/A sky130_fd_sc_hd__mux4_1
XFILLER_120_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23565_ _23577_/A _23565_/B vssd1 vssd1 vccd1 vccd1 _23566_/A sky130_fd_sc_hd__and2_1
X_26353_ _20547_/X _26353_/D vssd1 vssd1 vccd1 vccd1 _26353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20777_ _20853_/A vssd1 vssd1 vccd1 vccd1 _20777_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22516_ _22516_/A vssd1 vssd1 vccd1 vccd1 _22516_/X sky130_fd_sc_hd__clkbuf_1
X_25304_ _25304_/A _25304_/B vssd1 vssd1 vccd1 vccd1 _25329_/B sky130_fd_sc_hd__nand2_1
X_26284_ _20301_/X _26284_/D vssd1 vssd1 vccd1 vccd1 _26284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23496_ input30/X _23429_/A _23495_/X _23487_/X vssd1 vssd1 vccd1 vccd1 _27191_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_28023_ _28023_/A _15978_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_22447_ _22433_/X _22434_/X _22435_/X _22436_/X _22438_/X _22440_/X vssd1 vssd1 vccd1
+ vccd1 _22448_/A sky130_fd_sc_hd__mux4_1
X_25235_ _25250_/A _25235_/B vssd1 vssd1 vccd1 vccd1 _25242_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25166_ _25182_/A _25166_/B vssd1 vssd1 vccd1 vccd1 _25166_/Y sky130_fd_sc_hd__nand2_1
X_13180_ _27044_/Q _13179_/X _13199_/S vssd1 vssd1 vccd1 vccd1 _13181_/A sky130_fd_sc_hd__mux2_1
X_22378_ _22378_/A vssd1 vssd1 vccd1 vccd1 _22378_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24117_ _27406_/Q _24117_/B vssd1 vssd1 vccd1 vccd1 _24118_/A sky130_fd_sc_hd__and2_1
X_21329_ _21377_/A vssd1 vssd1 vccd1 vccd1 _21329_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25097_ _27977_/A _25096_/X _25104_/S vssd1 vssd1 vccd1 vccd1 _25098_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24048_ _27097_/Q _23860_/A _23861_/A _27129_/Q _23862_/A vssd1 vssd1 vccd1 vccd1
+ _24048_/X sky130_fd_sc_hd__a221o_1
XFILLER_81_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _16640_/A _16867_/X _16869_/Y vssd1 vssd1 vccd1 vccd1 _25615_/A sky130_fd_sc_hd__o21a_1
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27807_ _25680_/X _27807_/D vssd1 vssd1 vccd1 vccd1 _27807_/Q sky130_fd_sc_hd__dfxtp_1
X_15821_ _13150_/X _26089_/Q _15827_/S vssd1 vssd1 vccd1 vccd1 _15822_/A sky130_fd_sc_hd__mux2_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25999_ _26030_/CLK _25999_/D vssd1 vssd1 vccd1 vccd1 _25999_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18540_ _26295_/Q _26263_/Q _26231_/Q _26199_/Q _18458_/X _18481_/X vssd1 vssd1 vccd1
+ vccd1 _18540_/X sky130_fd_sc_hd__mux4_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _26118_/Q _15747_/X _15740_/X _15751_/Y vssd1 vssd1 vccd1 vccd1 _26118_/D
+ sky130_fd_sc_hd__a31o_1
X_27738_ _27748_/CLK _27738_/D vssd1 vssd1 vccd1 vccd1 _27738_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _12964_/A vssd1 vssd1 vccd1 vccd1 _27815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _15777_/A _14707_/B vssd1 vssd1 vccd1 vccd1 _14703_/Y sky130_fd_sc_hd__nor2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _18469_/X _18470_/X _18532_/S vssd1 vssd1 vccd1 vccd1 _18471_/X sky130_fd_sc_hd__mux2_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27669_ _27669_/CLK _27669_/D vssd1 vssd1 vccd1 vccd1 _27669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15683_ _13210_/X _26143_/Q _15689_/S vssd1 vssd1 vccd1 vccd1 _15684_/A sky130_fd_sc_hd__mux2_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_330 _25808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_341 _13334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_352 _14515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17422_ _23109_/A _27378_/Q _17674_/C vssd1 vssd1 vccd1 vccd1 _17601_/C sky130_fd_sc_hd__or3_1
XFILLER_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14634_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14646_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_363 _27593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_374 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17353_ _17303_/X _17352_/X _17342_/X vssd1 vssd1 vccd1 vccd1 _17353_/X sky130_fd_sc_hd__a21bo_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _26608_/Q _14563_/X _14553_/X _14564_/Y vssd1 vssd1 vccd1 vccd1 _26608_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _16304_/A _16304_/B vssd1 vssd1 vccd1 vccd1 _16304_/Y sky130_fd_sc_hd__nor2_1
X_13516_ _14482_/A vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__clkbuf_2
X_17284_ _27088_/Q _27120_/Q _17295_/S vssd1 vssd1 vccd1 vccd1 _17284_/X sky130_fd_sc_hd__mux2_1
X_14496_ _14530_/A vssd1 vssd1 vccd1 vccd1 _14496_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19023_ _19393_/A vssd1 vssd1 vccd1 vccd1 _19023_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16235_ _16235_/A _16235_/B _16235_/C vssd1 vssd1 vccd1 vccd1 _16235_/X sky130_fd_sc_hd__and3_1
X_13447_ _13546_/A vssd1 vssd1 vccd1 vccd1 _13471_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13378_ _13378_/A vssd1 vssd1 vccd1 vccd1 _26984_/D sky130_fd_sc_hd__clkbuf_1
X_16166_ _26052_/Q _16249_/B _16233_/C vssd1 vssd1 vccd1 vccd1 _16166_/X sky130_fd_sc_hd__and3_1
XFILLER_182_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15117_ _15117_/A vssd1 vssd1 vccd1 vccd1 _26394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _16374_/A vssd1 vssd1 vccd1 vccd1 _16098_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19925_ _25659_/A vssd1 vssd1 vccd1 vccd1 _20272_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15048_ _15116_/S vssd1 vssd1 vccd1 vccd1 _15057_/S sky130_fd_sc_hd__buf_2
XFILLER_102_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19856_ _19850_/X _19851_/X _19852_/X _19853_/X _19854_/X _19855_/X vssd1 vssd1 vccd1
+ vccd1 _19857_/A sky130_fd_sc_hd__mux4_1
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18807_ _19165_/A vssd1 vssd1 vccd1 vccd1 _18807_/X sky130_fd_sc_hd__clkbuf_4
X_19787_ _19787_/A vssd1 vssd1 vccd1 vccd1 _19787_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16999_ _17325_/A vssd1 vssd1 vccd1 vccd1 _17061_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18738_ _26030_/Q _17740_/X _18746_/S vssd1 vssd1 vccd1 vccd1 _18739_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18669_ _18669_/A vssd1 vssd1 vccd1 vccd1 _25999_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20700_ _20684_/X _20685_/X _20686_/X _20687_/X _20689_/X _20691_/X vssd1 vssd1 vccd1
+ vccd1 _20701_/A sky130_fd_sc_hd__mux4_1
XFILLER_52_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21680_ _21680_/A vssd1 vssd1 vccd1 vccd1 _21680_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20631_ _20631_/A vssd1 vssd1 vccd1 vccd1 _20631_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23350_ _27758_/Q vssd1 vssd1 vccd1 vccd1 _24844_/A sky130_fd_sc_hd__clkbuf_4
X_20562_ _20550_/X _20551_/X _20552_/X _20553_/X _20554_/X _20555_/X vssd1 vssd1 vccd1
+ vccd1 _20563_/A sky130_fd_sc_hd__mux4_1
XFILLER_177_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22301_ _22349_/A vssd1 vssd1 vccd1 vccd1 _22301_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23281_ input63/X vssd1 vssd1 vccd1 vccd1 _23281_/Y sky130_fd_sc_hd__inv_2
X_20493_ _20493_/A vssd1 vssd1 vccd1 vccd1 _20493_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25020_ _25917_/Q _25983_/Q _25816_/Q _26015_/Q _25009_/X _24983_/X vssd1 vssd1 vccd1
+ vccd1 _25020_/X sky130_fd_sc_hd__mux4_1
X_22232_ _22264_/A vssd1 vssd1 vccd1 vccd1 _22232_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22163_ _22157_/X _22158_/X _22159_/X _22160_/X _22161_/X _22162_/X vssd1 vssd1 vccd1
+ vccd1 _22164_/A sky130_fd_sc_hd__mux4_1
XFILLER_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21114_ _21114_/A vssd1 vssd1 vccd1 vccd1 _21114_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22094_ _22094_/A vssd1 vssd1 vccd1 vccd1 _22094_/X sky130_fd_sc_hd__clkbuf_1
X_26971_ _22708_/X _26971_/D vssd1 vssd1 vccd1 vccd1 _26971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25922_ _26020_/CLK _25922_/D vssd1 vssd1 vccd1 vccd1 _25922_/Q sky130_fd_sc_hd__dfxtp_1
X_21045_ _21217_/A vssd1 vssd1 vccd1 vccd1 _21114_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25853_ _27837_/CLK _25853_/D vssd1 vssd1 vccd1 vccd1 _25853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24804_ _24804_/A _24815_/B vssd1 vssd1 vccd1 vccd1 _24804_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25784_ _17492_/X _27847_/Q _25790_/S vssd1 vssd1 vccd1 vccd1 _25785_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22996_ _25638_/A vssd1 vssd1 vccd1 vccd1 _22996_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27523_ _27523_/CLK _27523_/D vssd1 vssd1 vccd1 vccd1 _27523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24735_ _24748_/A vssd1 vssd1 vccd1 vccd1 _24803_/A sky130_fd_sc_hd__clkbuf_2
X_21947_ _21930_/X _21932_/X _21934_/X _21936_/X _21937_/X _21938_/X vssd1 vssd1 vccd1
+ vccd1 _21948_/A sky130_fd_sc_hd__mux4_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27454_ _27454_/CLK _27454_/D vssd1 vssd1 vccd1 vccd1 _27454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21878_ _21878_/A vssd1 vssd1 vccd1 vccd1 _21878_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24666_ _24633_/A _24660_/X _24665_/X _24663_/X vssd1 vssd1 vccd1 vccd1 _27584_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26405_ _20729_/X _26405_/D vssd1 vssd1 vccd1 vccd1 _26405_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20829_ _20829_/A vssd1 vssd1 vccd1 vccd1 _20829_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23617_ _23617_/A _23617_/B vssd1 vssd1 vccd1 vccd1 _23618_/A sky130_fd_sc_hd__and2_1
X_27385_ _27386_/CLK _27385_/D vssd1 vssd1 vccd1 vccd1 _27385_/Q sky130_fd_sc_hd__dfxtp_1
X_24597_ _24597_/A vssd1 vssd1 vccd1 vccd1 _27558_/D sky130_fd_sc_hd__clkbuf_1
X_14350_ _14350_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _14350_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26336_ _20489_/X _26336_/D vssd1 vssd1 vccd1 vccd1 _26336_/Q sky130_fd_sc_hd__dfxtp_1
X_23548_ _23560_/A _23548_/B vssd1 vssd1 vccd1 vccd1 _23549_/A sky130_fd_sc_hd__and2_1
X_13301_ _13301_/A vssd1 vssd1 vccd1 vccd1 _27010_/D sky130_fd_sc_hd__clkbuf_1
X_14281_ _14369_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14281_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23479_ input23/X _23469_/X _23478_/X _23474_/X vssd1 vssd1 vccd1 vccd1 _27184_/D
+ sky130_fd_sc_hd__o211a_1
X_26267_ _20243_/X _26267_/D vssd1 vssd1 vccd1 vccd1 _26267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_28006_ _28006_/A _15860_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_16020_ _27481_/Q _27479_/Q _16020_/C vssd1 vssd1 vccd1 vccd1 _16020_/X sky130_fd_sc_hd__or3_1
X_13232_ _27336_/Q _13193_/A _13194_/A _27304_/Q _13231_/X vssd1 vssd1 vccd1 vccd1
+ _16177_/A sky130_fd_sc_hd__a221o_1
XFILLER_137_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25218_ _25218_/A _25218_/B vssd1 vssd1 vccd1 vccd1 _25220_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26198_ _20005_/X _26198_/D vssd1 vssd1 vccd1 vccd1 _26198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _13163_/A vssd1 vssd1 vccd1 vccd1 _27047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25149_ _25149_/A _25149_/B vssd1 vssd1 vccd1 vccd1 _25150_/B sky130_fd_sc_hd__nand2_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13094_ _14731_/A vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__buf_2
X_17971_ _17971_/A vssd1 vssd1 vccd1 vccd1 _25948_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19710_ _19726_/A vssd1 vssd1 vccd1 vccd1 _19710_/X sky130_fd_sc_hd__clkbuf_1
X_16922_ _27688_/Q vssd1 vssd1 vccd1 vccd1 _25108_/A sky130_fd_sc_hd__inv_2
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19641_ input4/X vssd1 vssd1 vccd1 vccd1 _22613_/A sky130_fd_sc_hd__buf_6
X_16853_ _16852_/A _16852_/B _16738_/A vssd1 vssd1 vccd1 vccd1 _16853_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15804_ _15804_/A vssd1 vssd1 vccd1 vccd1 _26097_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19572_ _19638_/A vssd1 vssd1 vccd1 vccd1 _19572_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16784_ _16733_/B _16708_/A _16774_/X _16774_/A _16711_/A vssd1 vssd1 vccd1 vccd1
+ _16785_/B sky130_fd_sc_hd__a32o_1
X_13996_ _14367_/A _14010_/B vssd1 vssd1 vccd1 vccd1 _13996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18523_ _26166_/Q _26102_/Q _27030_/Q _26998_/Q _17821_/X _17824_/X vssd1 vssd1 vccd1
+ vccd1 _18524_/A sky130_fd_sc_hd__mux4_1
X_15735_ _15761_/A vssd1 vssd1 vccd1 vccd1 _15745_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _12947_/A vssd1 vssd1 vccd1 vccd1 _27822_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _17995_/X _18449_/X _18451_/X _18453_/X _18352_/S vssd1 vssd1 vccd1 vccd1
+ _18466_/B sky130_fd_sc_hd__a221o_1
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15666_ _15666_/A vssd1 vssd1 vccd1 vccd1 _26151_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_160 _13382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _16298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_182 _14464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17405_ _19830_/A _19832_/A _19834_/A _19836_/A _19625_/A _19626_/A vssd1 vssd1 vccd1
+ vccd1 _17406_/A sky130_fd_sc_hd__mux4_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 _16243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ _26588_/Q _14615_/X _14605_/X _14616_/Y vssd1 vssd1 vccd1 vccd1 _26588_/D
+ sky130_fd_sc_hd__a31o_1
X_18385_ _18379_/X _18381_/X _18383_/X _18384_/X vssd1 vssd1 vccd1 vccd1 _18385_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15597_ _15608_/A vssd1 vssd1 vccd1 vccd1 _15606_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17336_ _17336_/A vssd1 vssd1 vccd1 vccd1 _27942_/A sky130_fd_sc_hd__clkbuf_1
X_14548_ _14548_/A vssd1 vssd1 vccd1 vccd1 _14602_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17267_ _25933_/Q _25999_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17268_/B sky130_fd_sc_hd__mux2_1
X_14479_ _16451_/A vssd1 vssd1 vccd1 vccd1 _15743_/A sky130_fd_sc_hd__buf_2
X_19006_ _18954_/X _19005_/X _18958_/X vssd1 vssd1 vccd1 vccd1 _19006_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16218_ _16218_/A _16221_/B _16235_/C vssd1 vssd1 vccd1 vccd1 _16218_/X sky130_fd_sc_hd__and3_1
XFILLER_174_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17198_ _27081_/Q _27113_/Q _17234_/S vssd1 vssd1 vccd1 vccd1 _17198_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16149_ _27399_/Q _16297_/B vssd1 vssd1 vccd1 vccd1 _16149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19908_ _19898_/X _19899_/X _19900_/X _19901_/X _19903_/X _19905_/X vssd1 vssd1 vccd1
+ vccd1 _19909_/A sky130_fd_sc_hd__mux4_1
XFILLER_69_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19839_ _19887_/A vssd1 vssd1 vccd1 vccd1 _19839_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22850_ _22850_/A vssd1 vssd1 vccd1 vccd1 _22850_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21801_ _21793_/X _21794_/X _21795_/X _21796_/X _21797_/X _21798_/X vssd1 vssd1 vccd1
+ vccd1 _21802_/A sky130_fd_sc_hd__mux4_1
X_22781_ _22767_/X _22768_/X _22769_/X _22770_/X _22771_/X _22772_/X vssd1 vssd1 vccd1
+ vccd1 _22782_/A sky130_fd_sc_hd__mux4_1
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21732_ _21732_/A vssd1 vssd1 vccd1 vccd1 _21732_/X sky130_fd_sc_hd__clkbuf_1
X_24520_ _24520_/A vssd1 vssd1 vccd1 vccd1 _27529_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21663_ _21647_/X _21648_/X _21649_/X _21650_/X _21652_/X _21654_/X vssd1 vssd1 vccd1
+ vccd1 _21664_/A sky130_fd_sc_hd__mux4_1
X_24451_ _24451_/A vssd1 vssd1 vccd1 vccd1 _27502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20614_ _20598_/X _20599_/X _20600_/X _20601_/X _20603_/X _20605_/X vssd1 vssd1 vccd1
+ vccd1 _20615_/A sky130_fd_sc_hd__mux4_1
X_23402_ _24823_/A _27233_/Q _27236_/Q _24737_/A vssd1 vssd1 vccd1 vccd1 _23402_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24382_ _25584_/A vssd1 vssd1 vccd1 vccd1 _25524_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_27170_ _27585_/CLK _27170_/D vssd1 vssd1 vccd1 vccd1 _27170_/Q sky130_fd_sc_hd__dfxtp_1
X_21594_ _21594_/A vssd1 vssd1 vccd1 vccd1 _21594_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26121_ _19737_/X _26121_/D vssd1 vssd1 vccd1 vccd1 _26121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23333_ _27262_/Q vssd1 vssd1 vccd1 vccd1 _23333_/Y sky130_fd_sc_hd__inv_2
X_20545_ _20545_/A vssd1 vssd1 vccd1 vccd1 _20545_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23264_ input59/X _23262_/Y _23263_/Y _27740_/Q vssd1 vssd1 vccd1 vccd1 _23264_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_26052_ _27333_/CLK _26052_/D vssd1 vssd1 vccd1 vccd1 _26052_/Q sky130_fd_sc_hd__dfxtp_1
X_20476_ _20464_/X _20465_/X _20466_/X _20467_/X _20468_/X _20469_/X vssd1 vssd1 vccd1
+ vccd1 _20477_/A sky130_fd_sc_hd__mux4_1
XFILLER_134_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22215_ _22263_/A vssd1 vssd1 vccd1 vccd1 _22215_/X sky130_fd_sc_hd__clkbuf_1
X_25003_ _25001_/X _25002_/X _25003_/S vssd1 vssd1 vccd1 vccd1 _25003_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23195_ _23252_/S vssd1 vssd1 vccd1 vccd1 _23204_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_134_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22146_ _22162_/A vssd1 vssd1 vccd1 vccd1 _22146_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22077_ _22067_/X _22068_/X _22069_/X _22070_/X _22071_/X _22072_/X vssd1 vssd1 vccd1
+ vccd1 _22078_/A sky130_fd_sc_hd__mux4_1
X_26954_ _22648_/X _26954_/D vssd1 vssd1 vccd1 vccd1 _26954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25905_ _26040_/CLK _25905_/D vssd1 vssd1 vccd1 vccd1 _25905_/Q sky130_fd_sc_hd__dfxtp_1
X_21028_ _21028_/A vssd1 vssd1 vccd1 vccd1 _21028_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26885_ _22408_/X _26885_/D vssd1 vssd1 vccd1 vccd1 _26885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25836_ _25900_/CLK _25836_/D vssd1 vssd1 vccd1 vccd1 _25836_/Q sky130_fd_sc_hd__dfxtp_1
X_13850_ _16014_/B vssd1 vssd1 vccd1 vccd1 _15695_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25767_ _25767_/A vssd1 vssd1 vccd1 vccd1 _27839_/D sky130_fd_sc_hd__clkbuf_1
X_13781_ _13874_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13781_/Y sky130_fd_sc_hd__nor2_1
X_22979_ _25659_/A vssd1 vssd1 vccd1 vccd1 _25638_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27506_ _27625_/CLK _27506_/D vssd1 vssd1 vccd1 vccd1 _27506_/Q sky130_fd_sc_hd__dfxtp_1
X_15520_ _15520_/A vssd1 vssd1 vccd1 vccd1 _26216_/D sky130_fd_sc_hd__clkbuf_1
X_24718_ _27603_/Q _24714_/X _24716_/X _24717_/X vssd1 vssd1 vccd1 vccd1 _27603_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25698_ _25698_/A vssd1 vssd1 vccd1 vccd1 _25698_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27437_ _27437_/CLK _27437_/D vssd1 vssd1 vccd1 vccd1 _27437_/Q sky130_fd_sc_hd__dfxtp_1
X_15451_ _26246_/Q _13382_/X _15451_/S vssd1 vssd1 vccd1 vccd1 _15452_/A sky130_fd_sc_hd__mux2_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24649_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24663_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _26655_/Q _14392_/X _14398_/X _14401_/Y vssd1 vssd1 vccd1 vccd1 _26655_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18170_ _18264_/A _18170_/B _18170_/C vssd1 vssd1 vccd1 vccd1 _18171_/A sky130_fd_sc_hd__and3_1
X_15382_ _14775_/X _26277_/Q _15390_/S vssd1 vssd1 vccd1 vccd1 _15383_/A sky130_fd_sc_hd__mux2_1
X_27368_ _27368_/CLK _27368_/D vssd1 vssd1 vccd1 vccd1 _27368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17121_ _25820_/Q _26019_/Q _17158_/S vssd1 vssd1 vccd1 vccd1 _17121_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14333_ _14333_/A _14335_/B vssd1 vssd1 vccd1 vccd1 _14333_/Y sky130_fd_sc_hd__nor2_1
X_26319_ _20423_/X _26319_/D vssd1 vssd1 vccd1 vccd1 _26319_/Q sky130_fd_sc_hd__dfxtp_1
X_27299_ _27299_/CLK _27299_/D vssd1 vssd1 vccd1 vccd1 _27299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17052_ _17116_/A vssd1 vssd1 vccd1 vccd1 _17052_/X sky130_fd_sc_hd__clkbuf_2
X_14264_ _26706_/Q _14256_/X _14258_/X _14263_/Y vssd1 vssd1 vccd1 vccd1 _26706_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16003_ _27483_/Q _27482_/Q _27480_/Q vssd1 vssd1 vccd1 vccd1 _16020_/C sky130_fd_sc_hd__or3_1
X_13215_ _16218_/A vssd1 vssd1 vccd1 vccd1 _14798_/A sky130_fd_sc_hd__buf_2
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _14372_/A _14200_/B vssd1 vssd1 vccd1 vccd1 _14195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13146_ _27050_/Q _13144_/X _13167_/S vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__mux2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17954_ _26814_/Q _26782_/Q _26750_/Q _26718_/Q _17863_/X _17890_/X vssd1 vssd1 vccd1
+ vccd1 _17954_/X sky130_fd_sc_hd__mux4_1
X_13077_ _13077_/A vssd1 vssd1 vccd1 vccd1 _14724_/A sky130_fd_sc_hd__clkbuf_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16905_ _16836_/A _16598_/A _16650_/A vssd1 vssd1 vccd1 vccd1 _16905_/X sky130_fd_sc_hd__o21ba_1
Xrepeater306 _27564_/CLK vssd1 vssd1 vccd1 vccd1 _27668_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater317 _27693_/CLK vssd1 vssd1 vccd1 vccd1 _27695_/CLK sky130_fd_sc_hd__clkbuf_1
X_17885_ _26940_/Q _26908_/Q _26876_/Q _26844_/Q _17789_/X _17791_/X vssd1 vssd1 vccd1
+ vccd1 _17885_/X sky130_fd_sc_hd__mux4_2
Xrepeater328 _27776_/CLK vssd1 vssd1 vccd1 vccd1 _27250_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater339 _27719_/CLK vssd1 vssd1 vccd1 vccd1 _27784_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16836_ _16836_/A vssd1 vssd1 vccd1 vccd1 _16836_/Y sky130_fd_sc_hd__inv_2
X_19624_ _19640_/A vssd1 vssd1 vccd1 vccd1 _19624_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19555_ _19555_/A _19555_/B vssd1 vssd1 vccd1 vccd1 _19555_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16767_ _16767_/A _16780_/B vssd1 vssd1 vccd1 vccd1 _16767_/Y sky130_fd_sc_hd__nand2_1
X_13979_ _26801_/Q _13969_/X _13965_/X _13978_/Y vssd1 vssd1 vccd1 vccd1 _26801_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18506_ _26421_/Q _26389_/Q _26357_/Q _26325_/Q _18462_/X _18486_/X vssd1 vssd1 vccd1
+ vccd1 _18506_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15718_ _15718_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19486_ _19486_/A vssd1 vssd1 vccd1 vccd1 _19486_/X sky130_fd_sc_hd__clkbuf_2
X_16698_ _16698_/A _16698_/B vssd1 vssd1 vccd1 vccd1 _16808_/B sky130_fd_sc_hd__and2_1
XFILLER_181_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18437_ _18437_/A vssd1 vssd1 vccd1 vccd1 _18437_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _15649_/A vssd1 vssd1 vccd1 vccd1 _26159_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18368_ _26159_/Q _26095_/Q _27023_/Q _26991_/Q _17821_/X _17824_/X vssd1 vssd1 vccd1
+ vccd1 _18369_/A sky130_fd_sc_hd__mux4_1
XFILLER_159_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ _17299_/X _17314_/X _17316_/X _17318_/X vssd1 vssd1 vccd1 vccd1 _17319_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_179_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18299_ _26156_/Q _26092_/Q _27020_/Q _26988_/Q _18298_/X _18228_/X vssd1 vssd1 vccd1
+ vccd1 _18300_/A sky130_fd_sc_hd__mux4_1
XFILLER_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20330_ _20318_/X _20319_/X _20320_/X _20321_/X _20322_/X _20323_/X vssd1 vssd1 vccd1
+ vccd1 _20331_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20261_ _20261_/A vssd1 vssd1 vccd1 vccd1 _20261_/X sky130_fd_sc_hd__clkbuf_1
X_22000_ _22000_/A vssd1 vssd1 vccd1 vccd1 _22000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_709 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20192_ _20181_/X _20183_/X _20185_/X _20187_/X _20188_/X _20189_/X vssd1 vssd1 vccd1
+ vccd1 _20193_/A sky130_fd_sc_hd__mux4_1
XFILLER_130_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23951_ _27086_/Q _27118_/Q _23986_/S vssd1 vssd1 vccd1 vccd1 _23951_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22902_ _22902_/A vssd1 vssd1 vccd1 vccd1 _22902_/X sky130_fd_sc_hd__clkbuf_1
X_26670_ _21656_/X _26670_/D vssd1 vssd1 vccd1 vccd1 _26670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23882_ _23929_/A vssd1 vssd1 vccd1 vccd1 _23882_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25621_ _23638_/B _27980_/A _25623_/S vssd1 vssd1 vccd1 vccd1 _25622_/A sky130_fd_sc_hd__mux2_1
X_22833_ _22821_/X _22822_/X _22823_/X _22824_/X _22825_/X _22826_/X vssd1 vssd1 vccd1
+ vccd1 _22834_/A sky130_fd_sc_hd__mux4_1
XFILLER_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25552_ _25552_/A vssd1 vssd1 vccd1 vccd1 _25552_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22764_ _22764_/A vssd1 vssd1 vccd1 vccd1 _22764_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24503_ _27588_/Q _24505_/B vssd1 vssd1 vccd1 vccd1 _24503_/X sky130_fd_sc_hd__or2_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21715_ _21705_/X _21706_/X _21707_/X _21708_/X _21709_/X _21710_/X vssd1 vssd1 vccd1
+ vccd1 _21716_/A sky130_fd_sc_hd__mux4_1
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22695_ _22681_/X _22682_/X _22683_/X _22684_/X _22685_/X _22686_/X vssd1 vssd1 vccd1
+ vccd1 _22696_/A sky130_fd_sc_hd__mux4_1
X_25483_ _25543_/A vssd1 vssd1 vccd1 vccd1 _25483_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27222_ _27222_/CLK _27222_/D vssd1 vssd1 vccd1 vccd1 _27222_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21646_ _21646_/A vssd1 vssd1 vccd1 vccd1 _21646_/X sky130_fd_sc_hd__clkbuf_1
X_24434_ _24434_/A vssd1 vssd1 vccd1 vccd1 _27495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27153_ _27153_/CLK _27153_/D vssd1 vssd1 vccd1 vccd1 _27153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21577_ _21561_/X _21562_/X _21563_/X _21564_/X _21566_/X _21568_/X vssd1 vssd1 vccd1
+ vccd1 _21578_/A sky130_fd_sc_hd__mux4_1
X_24365_ _24365_/A vssd1 vssd1 vccd1 vccd1 _27464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_60 _18268_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_71 _18442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_82 _18826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26104_ _19677_/X _26104_/D vssd1 vssd1 vccd1 vccd1 _26104_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_93 _19091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20528_ _20512_/X _20513_/X _20514_/X _20515_/X _20517_/X _20519_/X vssd1 vssd1 vccd1
+ vccd1 _20529_/A sky130_fd_sc_hd__mux4_1
X_23316_ _23257_/Y input52/X _23306_/Y input53/X vssd1 vssd1 vccd1 vccd1 _23316_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_165_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27084_ _27211_/CLK _27084_/D vssd1 vssd1 vccd1 vccd1 _27084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24296_ _16259_/Y _16260_/X _24269_/X vssd1 vssd1 vccd1 vccd1 _27427_/D sky130_fd_sc_hd__o21a_1
XFILLER_197_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26035_ _27092_/CLK _26035_/D vssd1 vssd1 vccd1 vccd1 _26035_/Q sky130_fd_sc_hd__dfxtp_1
X_23247_ _23247_/A vssd1 vssd1 vccd1 vccd1 _27158_/D sky130_fd_sc_hd__clkbuf_1
X_20459_ _20459_/A vssd1 vssd1 vccd1 vccd1 _20459_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13000_ _13000_/A vssd1 vssd1 vccd1 vccd1 _13009_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23178_ _27128_/Q _17772_/X _23180_/S vssd1 vssd1 vccd1 vccd1 _23179_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22129_ _22161_/A vssd1 vssd1 vccd1 vccd1 _22129_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27986_ _27986_/A _15986_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
XFILLER_153_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26937_ _22588_/X _26937_/D vssd1 vssd1 vccd1 vccd1 _26937_/Q sky130_fd_sc_hd__dfxtp_1
X_14951_ _14804_/X _26460_/Q _14951_/S vssd1 vssd1 vccd1 vccd1 _14952_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13902_ _13902_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13902_/Y sky130_fd_sc_hd__nor2_1
X_17670_ _17670_/A vssd1 vssd1 vccd1 vccd1 _25905_/D sky130_fd_sc_hd__clkbuf_1
X_26868_ _22344_/X _26868_/D vssd1 vssd1 vccd1 vccd1 _26868_/Q sky130_fd_sc_hd__dfxtp_1
X_14882_ _14882_/A vssd1 vssd1 vccd1 vccd1 _26491_/D sky130_fd_sc_hd__clkbuf_1
X_16621_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16621_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13833_ _13833_/A vssd1 vssd1 vccd1 vccd1 _13833_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25819_ _26018_/CLK _25819_/D vssd1 vssd1 vccd1 vccd1 _25819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26799_ _22100_/X _26799_/D vssd1 vssd1 vccd1 vccd1 _26799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19340_ _19409_/A _19340_/B vssd1 vssd1 vccd1 vccd1 _19340_/X sky130_fd_sc_hd__or2_1
X_16552_ _16826_/A _16552_/B vssd1 vssd1 vccd1 vccd1 _16552_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ _13847_/B vssd1 vssd1 vccd1 vccd1 _13764_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15503_ _15549_/S vssd1 vssd1 vccd1 vccd1 _15512_/S sky130_fd_sc_hd__buf_2
X_19271_ _26828_/Q _26796_/Q _26764_/Q _26732_/Q _19203_/X _19248_/X vssd1 vssd1 vccd1
+ vccd1 _19272_/B sky130_fd_sc_hd__mux4_1
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16483_ _16483_/A vssd1 vssd1 vccd1 vccd1 _16700_/A sky130_fd_sc_hd__clkbuf_2
X_13695_ _13876_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13695_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18222_ _18220_/X _18221_/X _18514_/S vssd1 vssd1 vccd1 vccd1 _18222_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15434_ _26254_/Q _13357_/X _15440_/S vssd1 vssd1 vccd1 vccd1 _15435_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ _18151_/X _18152_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18153_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_961 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15365_ _15365_/A vssd1 vssd1 vccd1 vccd1 _26285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ _17104_/A vssd1 vssd1 vccd1 vccd1 _27923_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14316_ _14403_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14316_/Y sky130_fd_sc_hd__nor2_1
X_18084_ _18084_/A _24392_/A vssd1 vssd1 vccd1 vccd1 _18084_/X sky130_fd_sc_hd__or2b_1
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15296_ _15296_/A vssd1 vssd1 vccd1 vccd1 _26315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17035_ _16985_/X _17028_/X _17031_/X _17034_/X vssd1 vssd1 vccd1 vccd1 _17035_/X
+ sky130_fd_sc_hd__o22a_1
X_14247_ _26712_/Q _14238_/X _14242_/X _14246_/Y vssd1 vssd1 vccd1 vccd1 _26712_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _26737_/Q _14173_/X _14167_/X _14177_/Y vssd1 vssd1 vccd1 vccd1 _26737_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13129_ _27053_/Q _13128_/X _13140_/S vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__mux2_1
XFILLER_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _18983_/X _18985_/X _19057_/S vssd1 vssd1 vccd1 vccd1 _18986_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater103 _27155_/CLK vssd1 vssd1 vccd1 vccd1 _27157_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_140_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater114 _27299_/CLK vssd1 vssd1 vccd1 vccd1 _27288_/CLK sky130_fd_sc_hd__clkbuf_1
X_17937_ _18324_/A vssd1 vssd1 vccd1 vccd1 _17937_/X sky130_fd_sc_hd__buf_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater125 _26037_/CLK vssd1 vssd1 vccd1 vccd1 _27149_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater136 _27094_/CLK vssd1 vssd1 vccd1 vccd1 _25996_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater147 _26040_/CLK vssd1 vssd1 vccd1 vccd1 _27160_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17868_ _17799_/X _17864_/X _17867_/X _24394_/A vssd1 vssd1 vccd1 vccd1 _17868_/X
+ sky130_fd_sc_hd__o211a_1
Xrepeater158 _25878_/CLK vssd1 vssd1 vccd1 vccd1 _27412_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater169 _27081_/CLK vssd1 vssd1 vccd1 vccd1 _25991_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19607_ _19639_/A vssd1 vssd1 vccd1 vccd1 _19607_/X sky130_fd_sc_hd__clkbuf_1
X_16819_ _16666_/Y _16665_/X _16818_/X vssd1 vssd1 vccd1 vccd1 _16819_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17799_ _18322_/A vssd1 vssd1 vccd1 vccd1 _17799_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19538_ _27823_/Q _26584_/Q _26456_/Q _26136_/Q _18829_/X _18831_/X vssd1 vssd1 vccd1
+ vccd1 _19538_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19469_ _19469_/A vssd1 vssd1 vccd1 vccd1 _19469_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21500_ _21564_/A vssd1 vssd1 vccd1 vccd1 _21500_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22480_ _22480_/A vssd1 vssd1 vccd1 vccd1 _22480_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21431_ _21463_/A vssd1 vssd1 vccd1 vccd1 _21431_/X sky130_fd_sc_hd__clkbuf_2
X_24150_ _24150_/A vssd1 vssd1 vccd1 vccd1 _27347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21362_ _21378_/A vssd1 vssd1 vccd1 vccd1 _21362_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23101_ _27094_/Q _17766_/X _23103_/S vssd1 vssd1 vccd1 vccd1 _23102_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20313_ _20313_/A vssd1 vssd1 vccd1 vccd1 _20313_/X sky130_fd_sc_hd__clkbuf_1
X_24081_ _24081_/A vssd1 vssd1 vccd1 vccd1 _27316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21293_ _21285_/X _21286_/X _21287_/X _21288_/X _21289_/X _21290_/X vssd1 vssd1 vccd1
+ vccd1 _21294_/A sky130_fd_sc_hd__mux4_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23032_ _23032_/A vssd1 vssd1 vccd1 vccd1 _23032_/X sky130_fd_sc_hd__clkbuf_1
X_20244_ _20232_/X _20233_/X _20234_/X _20235_/X _20236_/X _20237_/X vssd1 vssd1 vccd1
+ vccd1 _20245_/A sky130_fd_sc_hd__mux4_1
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27840_ _27840_/CLK _27840_/D vssd1 vssd1 vccd1 vccd1 _27840_/Q sky130_fd_sc_hd__dfxtp_1
X_20175_ _20175_/A vssd1 vssd1 vccd1 vccd1 _20175_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27771_ _27773_/CLK _27771_/D vssd1 vssd1 vccd1 vccd1 _27771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24983_ _25035_/A vssd1 vssd1 vccd1 vccd1 _24983_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26722_ _21838_/X _26722_/D vssd1 vssd1 vccd1 vccd1 _26722_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23934_ _27084_/Q _23907_/X _23908_/X _27116_/Q _23909_/X vssd1 vssd1 vccd1 vccd1
+ _23934_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26653_ _21596_/X _26653_/D vssd1 vssd1 vccd1 vccd1 _26653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23865_ _23849_/X _23859_/X _23863_/X _23864_/X vssd1 vssd1 vccd1 vccd1 _27281_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_199_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25604_ _18594_/A _25344_/B _25603_/X _25568_/A vssd1 vssd1 vccd1 vccd1 _25604_/X
+ sky130_fd_sc_hd__a211o_1
X_22816_ _22816_/A vssd1 vssd1 vccd1 vccd1 _22816_/X sky130_fd_sc_hd__clkbuf_1
X_26584_ _21356_/X _26584_/D vssd1 vssd1 vccd1 vccd1 _26584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23796_ _27070_/Q _27102_/Q _23796_/S vssd1 vssd1 vccd1 vccd1 _23796_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25535_ _27706_/Q _25509_/X _25510_/X vssd1 vssd1 vccd1 vccd1 _25535_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22747_ _22735_/X _22736_/X _22737_/X _22738_/X _22739_/X _22740_/X vssd1 vssd1 vccd1
+ vccd1 _22748_/A sky130_fd_sc_hd__mux4_1
XFILLER_77_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ _13884_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25466_ _25466_/A vssd1 vssd1 vccd1 vccd1 _25592_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22678_ _22678_/A vssd1 vssd1 vccd1 vccd1 _22678_/X sky130_fd_sc_hd__clkbuf_1
X_27205_ _27209_/CLK _27205_/D vssd1 vssd1 vccd1 vccd1 _27205_/Q sky130_fd_sc_hd__dfxtp_1
X_24417_ _24417_/A vssd1 vssd1 vccd1 vccd1 _27487_/D sky130_fd_sc_hd__clkbuf_1
X_21629_ _21615_/X _21616_/X _21617_/X _21618_/X _21619_/X _21620_/X vssd1 vssd1 vccd1
+ vccd1 _21630_/A sky130_fd_sc_hd__mux4_1
XFILLER_166_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25397_ _25397_/A vssd1 vssd1 vccd1 vccd1 _27737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15150_ _15150_/A vssd1 vssd1 vccd1 vccd1 _26380_/D sky130_fd_sc_hd__clkbuf_1
X_27136_ _27833_/CLK _27136_/D vssd1 vssd1 vccd1 vccd1 _27136_/Q sky130_fd_sc_hd__dfxtp_1
X_24348_ _27557_/Q _24350_/B vssd1 vssd1 vccd1 vccd1 _24349_/A sky130_fd_sc_hd__and2_1
XFILLER_166_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14101_ _14367_/A _14112_/B vssd1 vssd1 vccd1 vccd1 _14101_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15081_ _15103_/A vssd1 vssd1 vccd1 vccd1 _15090_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_10_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_856 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27067_ _27410_/CLK _27067_/D vssd1 vssd1 vccd1 vccd1 _27067_/Q sky130_fd_sc_hd__dfxtp_1
X_24279_ _24279_/A vssd1 vssd1 vccd1 vccd1 _24279_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14032_ _14032_/A vssd1 vssd1 vccd1 vccd1 _14047_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26018_ _26018_/CLK _26018_/D vssd1 vssd1 vccd1 vccd1 _26018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18840_ _19220_/A vssd1 vssd1 vccd1 vccd1 _18840_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18771_ _26810_/Q _26778_/Q _26746_/Q _26714_/Q _18767_/X _18770_/X vssd1 vssd1 vccd1
+ vccd1 _18772_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15983_ _15985_/A vssd1 vssd1 vccd1 vccd1 _15983_/Y sky130_fd_sc_hd__inv_2
X_27969_ _27969_/A _15868_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17722_ _25926_/Q _17721_/X _17722_/S vssd1 vssd1 vccd1 vccd1 _17723_/A sky130_fd_sc_hd__mux2_1
X_14934_ _14779_/X _26468_/Q _14940_/S vssd1 vssd1 vccd1 vccd1 _14935_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17653_ _17653_/A vssd1 vssd1 vccd1 vccd1 _25897_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14865_ _14865_/A vssd1 vssd1 vccd1 vccd1 _26499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16604_ _16604_/A _16604_/B vssd1 vssd1 vccd1 vccd1 _16604_/Y sky130_fd_sc_hd__xnor2_1
X_13816_ _26855_/Q _13806_/X _13807_/X _13815_/Y vssd1 vssd1 vccd1 vccd1 _26855_/D
+ sky130_fd_sc_hd__a31o_1
X_17584_ _17501_/X _25867_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17585_/A sky130_fd_sc_hd__mux2_1
X_14796_ _14795_/X _26527_/Q _14805_/S vssd1 vssd1 vccd1 vccd1 _14797_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19323_ _19320_/X _19322_/X _19346_/S vssd1 vssd1 vccd1 vccd1 _19323_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16535_ _16535_/A _16535_/B vssd1 vssd1 vccd1 vccd1 _16660_/A sky130_fd_sc_hd__xor2_1
X_13747_ _26880_/Q _13737_/X _13745_/X _13746_/Y vssd1 vssd1 vccd1 vccd1 _26880_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19254_ _26955_/Q _26923_/Q _26891_/Q _26859_/Q _19208_/X _19253_/X vssd1 vssd1 vccd1
+ vccd1 _19254_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ _16779_/B _16441_/B _16450_/A _16450_/B vssd1 vssd1 vccd1 vccd1 _16466_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_13678_ _13857_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13678_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18205_ _18150_/X _18197_/X _18204_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _18218_/B
+ sky130_fd_sc_hd__a211o_1
X_15417_ _15417_/A vssd1 vssd1 vccd1 vccd1 _26262_/D sky130_fd_sc_hd__clkbuf_1
X_19185_ _19182_/X _19184_/X _19211_/S vssd1 vssd1 vccd1 vccd1 _19185_/X sky130_fd_sc_hd__mux2_1
X_16397_ _16394_/X _16395_/Y _16737_/B _16396_/X vssd1 vssd1 vccd1 vccd1 _16397_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18136_ _17972_/X _18131_/X _18135_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _18146_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_106_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15348_ _15405_/S vssd1 vssd1 vccd1 vccd1 _15357_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_184_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18067_ _18067_/A _18066_/X vssd1 vssd1 vccd1 vccd1 _18067_/X sky130_fd_sc_hd__or2b_1
X_15279_ _15279_/A vssd1 vssd1 vccd1 vccd1 _26323_/D sky130_fd_sc_hd__clkbuf_1
X_17018_ _17266_/A vssd1 vssd1 vccd1 vccd1 _17071_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_99_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18969_ _18969_/A _18969_/B vssd1 vssd1 vccd1 vccd1 _18969_/X sky130_fd_sc_hd__or2_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21980_ _21980_/A vssd1 vssd1 vccd1 vccd1 _21980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20931_ _20921_/X _20922_/X _20923_/X _20924_/X _20925_/X _20926_/X vssd1 vssd1 vccd1
+ vccd1 _20932_/A sky130_fd_sc_hd__mux4_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20862_ _20848_/X _20849_/X _20850_/X _20851_/X _20852_/X _20853_/X vssd1 vssd1 vccd1
+ vccd1 _20863_/A sky130_fd_sc_hd__mux4_1
X_23650_ _23650_/A _23650_/B vssd1 vssd1 vccd1 vccd1 _23707_/A sky130_fd_sc_hd__nand2_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22601_ _22593_/X _22594_/X _22595_/X _22596_/X _22597_/X _22598_/X vssd1 vssd1 vccd1
+ vccd1 _22602_/A sky130_fd_sc_hd__mux4_1
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23581_ _27773_/Q _27215_/Q _23595_/S vssd1 vssd1 vccd1 vccd1 _23582_/B sky130_fd_sc_hd__mux2_1
X_20793_ _22540_/A vssd1 vssd1 vccd1 vccd1 _21145_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25320_ _25320_/A _25320_/B vssd1 vssd1 vccd1 vccd1 _25321_/B sky130_fd_sc_hd__or2_1
X_22532_ _22532_/A vssd1 vssd1 vccd1 vccd1 _22532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25251_ _25243_/B _25250_/X _25241_/B vssd1 vssd1 vccd1 vccd1 _25252_/B sky130_fd_sc_hd__o21a_1
X_22463_ _22452_/X _22454_/X _22456_/X _22458_/X _22459_/X _22460_/X vssd1 vssd1 vccd1
+ vccd1 _22464_/A sky130_fd_sc_hd__mux4_1
X_24202_ _27754_/Q vssd1 vssd1 vccd1 vccd1 _25733_/A sky130_fd_sc_hd__buf_2
XFILLER_185_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21414_ _21478_/A vssd1 vssd1 vccd1 vccd1 _21414_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22394_ _22394_/A vssd1 vssd1 vccd1 vccd1 _22394_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25182_ _25182_/A _25182_/B vssd1 vssd1 vccd1 vccd1 _25182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21345_ _21377_/A vssd1 vssd1 vccd1 vccd1 _21345_/X sky130_fd_sc_hd__clkbuf_2
X_24133_ _24133_/A vssd1 vssd1 vccd1 vccd1 _27339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21276_ _21276_/A vssd1 vssd1 vccd1 vccd1 _21276_/X sky130_fd_sc_hd__clkbuf_1
X_24064_ _27382_/Q _24072_/B vssd1 vssd1 vccd1 vccd1 _24065_/A sky130_fd_sc_hd__and2_1
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20227_ _20227_/A vssd1 vssd1 vccd1 vccd1 _20227_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23015_ _23009_/X _23010_/X _23011_/X _23012_/X _23013_/X _23014_/X vssd1 vssd1 vccd1
+ vccd1 _23016_/A sky130_fd_sc_hd__mux4_1
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27823_ _25730_/X _27823_/D vssd1 vssd1 vccd1 vccd1 _27823_/Q sky130_fd_sc_hd__dfxtp_1
X_20158_ _20146_/X _20147_/X _20148_/X _20149_/X _20150_/X _20151_/X vssd1 vssd1 vccd1
+ vccd1 _20159_/A sky130_fd_sc_hd__mux4_1
XFILLER_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27754_ _27754_/CLK _27754_/D vssd1 vssd1 vccd1 vccd1 _27754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ _12980_/A vssd1 vssd1 vccd1 vccd1 _27808_/D sky130_fd_sc_hd__clkbuf_1
X_24966_ _24969_/B _24966_/B vssd1 vssd1 vccd1 vccd1 _24967_/B sky130_fd_sc_hd__nand2_1
X_20089_ _20089_/A vssd1 vssd1 vccd1 vccd1 _20089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26705_ _21784_/X _26705_/D vssd1 vssd1 vccd1 vccd1 _26705_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23917_ _23915_/X _23916_/X _23940_/S vssd1 vssd1 vccd1 vccd1 _23917_/X sky130_fd_sc_hd__mux2_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27685_ _27686_/CLK _27685_/D vssd1 vssd1 vccd1 vccd1 _27976_/A sky130_fd_sc_hd__dfxtp_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24897_ _24893_/A _24896_/C _27769_/Q vssd1 vssd1 vccd1 vccd1 _24898_/B sky130_fd_sc_hd__a21oi_1
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26636_ _21538_/X _26636_/D vssd1 vssd1 vccd1 vccd1 _26636_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _26577_/Q _14645_/X _14640_/X _14649_/Y vssd1 vssd1 vccd1 vccd1 _26577_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23848_ _23800_/X _23846_/X _23847_/X _23816_/X vssd1 vssd1 vccd1 vccd1 _27280_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13601_ _26933_/Q _13599_/X _13587_/X _13600_/Y vssd1 vssd1 vccd1 vccd1 _26933_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14581_ _26602_/Q _14576_/X _14579_/X _14580_/Y vssd1 vssd1 vccd1 vccd1 _26602_/D
+ sky130_fd_sc_hd__a31o_1
X_26567_ _21296_/X _26567_/D vssd1 vssd1 vccd1 vccd1 _26567_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23779_ _25914_/Q _25980_/Q _25813_/Q _26012_/Q _23747_/X _23749_/X vssd1 vssd1 vccd1
+ vccd1 _23779_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16320_ _16598_/A _16598_/B vssd1 vssd1 vccd1 vccd1 _16902_/A sky130_fd_sc_hd__and2_1
X_13532_ _14493_/A vssd1 vssd1 vccd1 vccd1 _13913_/A sky130_fd_sc_hd__clkbuf_2
X_25518_ _25517_/X _25492_/X _25493_/X _24889_/B _25494_/X vssd1 vssd1 vccd1 vccd1
+ _25518_/X sky130_fd_sc_hd__o311a_1
XFILLER_129_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26498_ _21054_/X _26498_/D vssd1 vssd1 vccd1 vccd1 _26498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _24287_/A _27533_/Q _16254_/S vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__mux2_1
X_13463_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__clkbuf_2
X_25449_ _25569_/A vssd1 vssd1 vccd1 vccd1 _25449_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15202_ _15202_/A vssd1 vssd1 vccd1 vccd1 _26357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16182_ _16182_/A _16215_/B _16197_/C vssd1 vssd1 vccd1 vccd1 _16182_/X sky130_fd_sc_hd__and3_1
X_13394_ _13394_/A vssd1 vssd1 vccd1 vccd1 _26979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27119_ _27296_/CLK _27119_/D vssd1 vssd1 vccd1 vccd1 _27119_/Q sky130_fd_sc_hd__dfxtp_1
X_15133_ _15133_/A vssd1 vssd1 vccd1 vccd1 _26388_/D sky130_fd_sc_hd__clkbuf_1
X_27995__461 vssd1 vssd1 vccd1 vccd1 _27995__461/HI _27995_/A sky130_fd_sc_hd__conb_1
XFILLER_182_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19941_ _19989_/A vssd1 vssd1 vccd1 vccd1 _19941_/X sky130_fd_sc_hd__clkbuf_1
X_15064_ _14734_/X _26418_/Q _15068_/S vssd1 vssd1 vccd1 vccd1 _15065_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ _26791_/Q _14005_/X _14001_/X _14014_/Y vssd1 vssd1 vccd1 vccd1 _26791_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19872_ _19866_/X _19867_/X _19868_/X _19869_/X _19870_/X _19871_/X vssd1 vssd1 vccd1
+ vccd1 _19873_/A sky130_fd_sc_hd__mux4_1
X_18823_ _19297_/A vssd1 vssd1 vccd1 vccd1 _19343_/A sky130_fd_sc_hd__buf_4
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18754_ _18754_/A vssd1 vssd1 vccd1 vccd1 _26037_/D sky130_fd_sc_hd__clkbuf_1
X_15966_ _15967_/A vssd1 vssd1 vccd1 vccd1 _15966_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17705_ _27417_/Q vssd1 vssd1 vccd1 vccd1 _17705_/X sky130_fd_sc_hd__clkbuf_2
X_14917_ _14917_/A vssd1 vssd1 vccd1 vccd1 _26476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15897_ _15899_/A vssd1 vssd1 vccd1 vccd1 _15897_/Y sky130_fd_sc_hd__inv_2
X_18685_ _26007_/Q _17769_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _18686_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17636_ _17658_/A vssd1 vssd1 vccd1 vccd1 _17645_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14848_ _14870_/A vssd1 vssd1 vccd1 vccd1 _14857_/S sky130_fd_sc_hd__buf_2
XFILLER_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_527 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17567_ _17476_/X _25859_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17568_/A sky130_fd_sc_hd__mux2_1
X_14779_ _14779_/A vssd1 vssd1 vccd1 vccd1 _14779_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16518_ _16292_/B _16292_/C _16292_/D _16106_/A vssd1 vssd1 vccd1 vccd1 _16519_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_17_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19306_ _18929_/A _19305_/X _18932_/A vssd1 vssd1 vccd1 vccd1 _19306_/X sky130_fd_sc_hd__o21a_1
XFILLER_177_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _27431_/Q vssd1 vssd1 vccd1 vccd1 _17498_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19237_ _19261_/A _19237_/B vssd1 vssd1 vccd1 vccd1 _19237_/X sky130_fd_sc_hd__or2_1
X_16449_ _16767_/A _16449_/B vssd1 vssd1 vccd1 vccd1 _16450_/B sky130_fd_sc_hd__xnor2_2
XFILLER_104_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19168_ _26279_/Q _26247_/Q _26215_/Q _26183_/Q _19144_/X _19074_/X vssd1 vssd1 vccd1
+ vccd1 _19168_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18119_ _26404_/Q _26372_/Q _26340_/Q _26308_/Q _18048_/X _18073_/X vssd1 vssd1 vccd1
+ vccd1 _18119_/X sky130_fd_sc_hd__mux4_1
X_19099_ _19073_/X _19098_/X _19076_/X vssd1 vssd1 vccd1 vccd1 _19099_/X sky130_fd_sc_hd__o21a_1
XFILLER_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21130_ _21199_/A vssd1 vssd1 vccd1 vccd1 _21130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21061_ _21147_/A vssd1 vssd1 vccd1 vccd1 _21127_/A sky130_fd_sc_hd__buf_2
XFILLER_63_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20012_ _20270_/A vssd1 vssd1 vccd1 vccd1 _20078_/A sky130_fd_sc_hd__buf_2
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24820_ _24841_/A vssd1 vssd1 vccd1 vccd1 _25601_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24751_ _27614_/Q _24742_/X _24750_/Y _24746_/X vssd1 vssd1 vccd1 vccd1 _27614_/D
+ sky130_fd_sc_hd__o211a_1
X_21963_ _21949_/X _21950_/X _21951_/X _21952_/X _21953_/X _21954_/X vssd1 vssd1 vccd1
+ vccd1 _21964_/A sky130_fd_sc_hd__mux4_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23702_ _23702_/A vssd1 vssd1 vccd1 vccd1 _27255_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _20914_/A vssd1 vssd1 vccd1 vccd1 _20914_/X sky130_fd_sc_hd__clkbuf_1
X_27470_ _27473_/CLK _27470_/D vssd1 vssd1 vccd1 vccd1 _27470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24682_ _27590_/Q _24673_/X _24681_/X _24677_/X vssd1 vssd1 vccd1 vccd1 _27590_/D
+ sky130_fd_sc_hd__o211a_1
X_21894_ _21894_/A vssd1 vssd1 vccd1 vccd1 _21894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26421_ _20781_/X _26421_/D vssd1 vssd1 vccd1 vccd1 _26421_/Q sky130_fd_sc_hd__dfxtp_1
X_23633_ _25004_/S vssd1 vssd1 vccd1 vccd1 _23638_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20845_/A vssd1 vssd1 vccd1 vccd1 _20845_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26352_ _20545_/X _26352_/D vssd1 vssd1 vccd1 vccd1 _26352_/Q sky130_fd_sc_hd__dfxtp_1
X_23564_ _24893_/A _27210_/Q _23576_/S vssd1 vssd1 vccd1 vccd1 _23565_/B sky130_fd_sc_hd__mux2_1
XFILLER_167_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20776_ _20776_/A vssd1 vssd1 vccd1 vccd1 _20853_/A sky130_fd_sc_hd__buf_2
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25303_ _25310_/A _27511_/Q vssd1 vssd1 vccd1 vccd1 _25304_/B sky130_fd_sc_hd__nand2_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22515_ _22503_/X _22504_/X _22505_/X _22506_/X _22507_/X _22508_/X vssd1 vssd1 vccd1
+ vccd1 _22516_/A sky130_fd_sc_hd__mux4_1
XFILLER_195_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26283_ _20299_/X _26283_/D vssd1 vssd1 vccd1 vccd1 _26283_/Q sky130_fd_sc_hd__dfxtp_1
X_23495_ _27191_/Q _23495_/B vssd1 vssd1 vccd1 vccd1 _23495_/X sky130_fd_sc_hd__or2_1
XFILLER_202_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_28022_ _28022_/A _15979_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
X_25234_ _27535_/Q _27503_/Q vssd1 vssd1 vccd1 vccd1 _25235_/B sky130_fd_sc_hd__nor2_1
XFILLER_167_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22446_ _22446_/A vssd1 vssd1 vccd1 vccd1 _22446_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25165_ _25165_/A _25165_/B vssd1 vssd1 vccd1 vccd1 _25166_/B sky130_fd_sc_hd__xor2_1
X_22377_ _22366_/X _22368_/X _22370_/X _22372_/X _22373_/X _22374_/X vssd1 vssd1 vccd1
+ vccd1 _22378_/A sky130_fd_sc_hd__mux4_1
XFILLER_135_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24116_ _24116_/A vssd1 vssd1 vccd1 vccd1 _27332_/D sky130_fd_sc_hd__clkbuf_1
X_21328_ _21392_/A vssd1 vssd1 vccd1 vccd1 _21328_/X sky130_fd_sc_hd__clkbuf_1
X_25096_ _25094_/X _25095_/X _25103_/S vssd1 vssd1 vccd1 vccd1 _25096_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21259_ _21253_/X _21254_/X _21255_/X _21256_/X _21257_/X _21258_/X vssd1 vssd1 vccd1
+ vccd1 _21260_/A sky130_fd_sc_hd__mux4_1
X_24047_ _24045_/X _24046_/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24047_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_551 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15820_ _15820_/A vssd1 vssd1 vccd1 vccd1 _26090_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27806_ _25672_/X _27806_/D vssd1 vssd1 vccd1 vccd1 _27806_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25998_ _27121_/CLK _25998_/D vssd1 vssd1 vccd1 vccd1 _25998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15751_ _15751_/A _15758_/B vssd1 vssd1 vccd1 vccd1 _15751_/Y sky130_fd_sc_hd__nor2_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27737_ _27737_/CLK _27737_/D vssd1 vssd1 vccd1 vccd1 _27737_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24949_ _24962_/A _24949_/B vssd1 vssd1 vccd1 vccd1 _24949_/Y sky130_fd_sc_hd__nand2_1
X_12963_ _27815_/Q _12965_/B vssd1 vssd1 vccd1 vccd1 _12964_/A sky130_fd_sc_hd__and2_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _26557_/Q _14698_/X _14693_/X _14701_/Y vssd1 vssd1 vccd1 vccd1 _26557_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _26964_/Q _26932_/Q _26900_/Q _26868_/Q _18403_/X _18427_/X vssd1 vssd1 vccd1
+ vccd1 _18470_/X sky130_fd_sc_hd__mux4_1
X_27668_ _27668_/CLK _27668_/D vssd1 vssd1 vccd1 vccd1 _27668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15682_ _15682_/A vssd1 vssd1 vccd1 vccd1 _26144_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_320 _19045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 _13244_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _27375_/Q _24003_/A vssd1 vssd1 vccd1 vccd1 _17674_/C sky130_fd_sc_hd__nand2_1
XANTENNA_342 _13347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26619_ _21474_/X _26619_/D vssd1 vssd1 vccd1 vccd1 _26619_/Q sky130_fd_sc_hd__dfxtp_1
X_14633_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 _14527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27599_ _27602_/CLK _27599_/D vssd1 vssd1 vccd1 vccd1 _27599_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_364 _27601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _25839_/Q _26038_/Q _17382_/S vssd1 vssd1 vccd1 vccd1 _17352_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _15725_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14564_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16836_/A _16593_/B _16595_/B vssd1 vssd1 vccd1 vccd1 _16304_/B sky130_fd_sc_hd__and3_1
XFILLER_202_875 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ _27349_/Q _13450_/X _13451_/X _27317_/Q _13153_/X vssd1 vssd1 vccd1 vccd1
+ _14482_/A sky130_fd_sc_hd__a221oi_4
X_17283_ _17238_/X _17276_/X _17279_/X _17282_/X vssd1 vssd1 vccd1 vccd1 _17283_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14495_ _26629_/Q _14478_/X _14492_/X _14494_/Y vssd1 vssd1 vccd1 vccd1 _26629_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19022_ _19324_/A vssd1 vssd1 vccd1 vccd1 _19022_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16234_ _27385_/Q _16244_/B _16244_/C vssd1 vssd1 vccd1 vccd1 _16234_/X sky130_fd_sc_hd__and3_1
XFILLER_174_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ _13456_/A vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_186_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16165_ _16108_/A _16445_/A _16162_/Y _16445_/B _16164_/X vssd1 vssd1 vccd1 vccd1
+ _16422_/A sky130_fd_sc_hd__o41a_1
XFILLER_177_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13377_ _26984_/Q _13376_/X _13383_/S vssd1 vssd1 vccd1 vccd1 _13378_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15116_ _14810_/X _26394_/Q _15116_/S vssd1 vssd1 vccd1 vccd1 _15117_/A sky130_fd_sc_hd__mux2_1
X_16096_ _16310_/A vssd1 vssd1 vccd1 vccd1 _16374_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19924_ _19990_/A vssd1 vssd1 vccd1 vccd1 _19924_/X sky130_fd_sc_hd__clkbuf_1
X_15047_ _15103_/A vssd1 vssd1 vccd1 vccd1 _15116_/S sky130_fd_sc_hd__buf_2
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19855_ _19887_/A vssd1 vssd1 vccd1 vccd1 _19855_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18806_ _27599_/Q vssd1 vssd1 vccd1 vccd1 _19165_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19786_ _19780_/X _19781_/X _19782_/X _19783_/X _19784_/X _19785_/X vssd1 vssd1 vccd1
+ vccd1 _19787_/A sky130_fd_sc_hd__mux4_1
XFILLER_37_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16998_ _17303_/A vssd1 vssd1 vccd1 vccd1 _16998_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18737_ _18748_/A vssd1 vssd1 vccd1 vccd1 _18746_/S sky130_fd_sc_hd__clkbuf_2
X_15949_ _15949_/A vssd1 vssd1 vccd1 vccd1 _15949_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18668_ _25999_/Q _17744_/X _18674_/S vssd1 vssd1 vccd1 vccd1 _18669_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17619_ _17447_/X _25882_/Q _17623_/S vssd1 vssd1 vccd1 vccd1 _17620_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18599_ _25568_/A _25113_/A vssd1 vssd1 vccd1 vccd1 _18599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20630_ _20617_/X _20619_/X _20621_/X _20623_/X _20624_/X _20625_/X vssd1 vssd1 vccd1
+ vccd1 _20631_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20561_ _20561_/A vssd1 vssd1 vccd1 vccd1 _20561_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22300_ _22348_/A vssd1 vssd1 vccd1 vccd1 _22300_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20492_ _20480_/X _20481_/X _20482_/X _20483_/X _20484_/X _20485_/X vssd1 vssd1 vccd1
+ vccd1 _20493_/A sky130_fd_sc_hd__mux4_1
X_23280_ _27721_/Q vssd1 vssd1 vccd1 vccd1 _23280_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22231_ _22263_/A vssd1 vssd1 vccd1 vccd1 _22231_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22162_ _22162_/A vssd1 vssd1 vccd1 vccd1 _22162_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21113_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22093_ _22083_/X _22084_/X _22085_/X _22086_/X _22088_/X _22090_/X vssd1 vssd1 vccd1
+ vccd1 _22094_/A sky130_fd_sc_hd__mux4_1
X_26970_ _22706_/X _26970_/D vssd1 vssd1 vccd1 vccd1 _26970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25921_ _25987_/CLK _25921_/D vssd1 vssd1 vccd1 vccd1 _25921_/Q sky130_fd_sc_hd__dfxtp_1
X_21044_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25852_ _27140_/CLK _25852_/D vssd1 vssd1 vccd1 vccd1 _25852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24803_ _24803_/A vssd1 vssd1 vccd1 vccd1 _24815_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25783_ _25783_/A vssd1 vssd1 vccd1 vccd1 _27846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22995_ _25637_/A vssd1 vssd1 vccd1 vccd1 _22995_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27522_ _27523_/CLK _27522_/D vssd1 vssd1 vccd1 vccd1 _27522_/Q sky130_fd_sc_hd__dfxtp_1
X_24734_ _27610_/Q _24727_/X _24733_/Y _24729_/X vssd1 vssd1 vccd1 vccd1 _27610_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21946_ _21946_/A vssd1 vssd1 vccd1 vccd1 _21946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_972 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27453_ _27454_/CLK _27453_/D vssd1 vssd1 vccd1 vccd1 _27453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24665_ _27168_/Q _24671_/B vssd1 vssd1 vccd1 vccd1 _24665_/X sky130_fd_sc_hd__or2_1
X_21877_ _21863_/X _21864_/X _21865_/X _21866_/X _21867_/X _21868_/X vssd1 vssd1 vccd1
+ vccd1 _21878_/A sky130_fd_sc_hd__mux4_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26404_ _20721_/X _26404_/D vssd1 vssd1 vccd1 vccd1 _26404_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23616_ _24960_/A _27224_/Q _23616_/S vssd1 vssd1 vccd1 vccd1 _23617_/B sky130_fd_sc_hd__mux2_1
X_20828_ _20816_/X _20817_/X _20818_/X _20819_/X _20820_/X _20821_/X vssd1 vssd1 vccd1
+ vccd1 _20829_/A sky130_fd_sc_hd__mux4_1
X_27384_ _27386_/CLK _27384_/D vssd1 vssd1 vccd1 vccd1 _27384_/Q sky130_fd_sc_hd__dfxtp_1
X_24596_ _27658_/Q _24598_/B vssd1 vssd1 vccd1 vccd1 _24597_/A sky130_fd_sc_hd__and2_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26335_ _20487_/X _26335_/D vssd1 vssd1 vccd1 vccd1 _26335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23547_ _27763_/Q _27205_/Q _23559_/S vssd1 vssd1 vccd1 vccd1 _23548_/B sky130_fd_sc_hd__mux2_1
X_20759_ _20759_/A vssd1 vssd1 vccd1 vccd1 _20759_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13300_ _27010_/Q _13190_/X _13302_/S vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__mux2_1
XFILLER_195_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14280_ _26700_/Q _14270_/X _14271_/X _14279_/Y vssd1 vssd1 vccd1 vccd1 _26700_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_183_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26266_ _20241_/X _26266_/D vssd1 vssd1 vccd1 vccd1 _26266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23478_ _27184_/Q _23483_/B vssd1 vssd1 vccd1 vccd1 _23478_/X sky130_fd_sc_hd__or2_1
X_28005_ _28005_/A _15861_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_25217_ _27533_/Q _27501_/Q vssd1 vssd1 vccd1 vccd1 _25218_/B sky130_fd_sc_hd__or2_1
X_13231_ _27272_/Q _13231_/B vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__and2_2
XFILLER_183_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22429_ _22417_/X _22418_/X _22419_/X _22420_/X _22421_/X _22422_/X vssd1 vssd1 vccd1
+ vccd1 _22430_/A sky130_fd_sc_hd__mux4_1
X_26197_ _20003_/X _26197_/D vssd1 vssd1 vccd1 vccd1 _26197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25148_ _25129_/A _25126_/X _25129_/B _25136_/A _25127_/A vssd1 vssd1 vccd1 vccd1
+ _25149_/B sky130_fd_sc_hd__a311o_1
X_13162_ _27047_/Q _13161_/X _13167_/S vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25079_ _25924_/Q _25990_/Q _25823_/Q _26022_/Q _25052_/X _25070_/X vssd1 vssd1 vccd1
+ vccd1 _25079_/X sky130_fd_sc_hd__mux4_1
X_17970_ _18028_/A _17970_/B _17970_/C vssd1 vssd1 vccd1 vccd1 _17971_/A sky130_fd_sc_hd__and3_1
X_13093_ _27360_/Q _13090_/X _13091_/X _27328_/Q _13092_/X vssd1 vssd1 vccd1 vccd1
+ _14731_/A sky130_fd_sc_hd__a221o_2
XFILLER_3_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16921_ _27574_/Q vssd1 vssd1 vccd1 vccd1 _25584_/A sky130_fd_sc_hd__inv_2
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19640_ _19640_/A vssd1 vssd1 vccd1 vccd1 _19640_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16852_ _16852_/A _16852_/B vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15803_ _13105_/X _26097_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15804_/A sky130_fd_sc_hd__mux2_1
X_19571_ _19832_/A vssd1 vssd1 vccd1 vccd1 _19638_/A sky130_fd_sc_hd__clkbuf_2
X_16783_ _16783_/A vssd1 vssd1 vccd1 vccd1 _16783_/Y sky130_fd_sc_hd__inv_2
X_13995_ _14032_/A vssd1 vssd1 vccd1 vccd1 _14010_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15734_ _24980_/S vssd1 vssd1 vccd1 vccd1 _15734_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18522_ _18520_/X _18521_/X _18522_/S vssd1 vssd1 vccd1 vccd1 _18522_/X sky130_fd_sc_hd__mux2_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _27822_/Q _12952_/B vssd1 vssd1 vccd1 vccd1 _12947_/A sky130_fd_sc_hd__and2_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _17912_/X _18452_/X _17915_/X vssd1 vssd1 vccd1 vccd1 _18453_/X sky130_fd_sc_hd__o21a_1
X_15665_ _13161_/X _26151_/Q _15667_/S vssd1 vssd1 vccd1 vccd1 _15666_/A sky130_fd_sc_hd__mux2_1
XFILLER_179_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_150 _13184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _16298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14616_ _15777_/A _14620_/B vssd1 vssd1 vccd1 vccd1 _14616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17404_ _25641_/A vssd1 vssd1 vccd1 vccd1 _19626_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _16277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18384_ _18384_/A vssd1 vssd1 vccd1 vccd1 _18384_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_194 _16243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15596_ _15596_/A vssd1 vssd1 vccd1 vccd1 _26182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _27221_/Q _17334_/X _17367_/S vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14547_ _26614_/Q _14530_/X _14536_/X _14546_/Y vssd1 vssd1 vccd1 vccd1 _26614_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_418 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17266_ _17266_/A vssd1 vssd1 vccd1 vccd1 _17315_/S sky130_fd_sc_hd__buf_2
X_14478_ _14530_/A vssd1 vssd1 vccd1 vccd1 _14478_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_186_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19005_ _26272_/Q _26240_/Q _26208_/Q _26176_/Q _18859_/X _18955_/X vssd1 vssd1 vccd1
+ vccd1 _19005_/X sky130_fd_sc_hd__mux4_1
X_16217_ _17674_/B _16233_/B vssd1 vssd1 vccd1 vccd1 _16217_/Y sky130_fd_sc_hd__nor2_1
X_13429_ _13583_/B vssd1 vssd1 vccd1 vccd1 _13429_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17197_ _17177_/X _17192_/X _17194_/X _17196_/X vssd1 vssd1 vccd1 vccd1 _17197_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16148_ _26065_/Q vssd1 vssd1 vccd1 vccd1 _16148_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _16648_/A vssd1 vssd1 vccd1 vccd1 _16559_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19907_ _19907_/A vssd1 vssd1 vccd1 vccd1 _19907_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19838_ _19886_/A vssd1 vssd1 vccd1 vccd1 _19838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_574 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
X_19769_ _19801_/A vssd1 vssd1 vccd1 vccd1 _19769_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21800_ _21800_/A vssd1 vssd1 vccd1 vccd1 _21800_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22780_ _22780_/A vssd1 vssd1 vccd1 vccd1 _22780_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21731_ _21721_/X _21722_/X _21723_/X _21724_/X _21725_/X _21726_/X vssd1 vssd1 vccd1
+ vccd1 _21732_/A sky130_fd_sc_hd__mux4_1
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24450_ _27623_/Q _24456_/B vssd1 vssd1 vccd1 vccd1 _24451_/A sky130_fd_sc_hd__and2_1
X_21662_ _21662_/A vssd1 vssd1 vccd1 vccd1 _21662_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23401_ _27756_/Q vssd1 vssd1 vccd1 vccd1 _24737_/A sky130_fd_sc_hd__inv_2
XFILLER_178_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20613_ _20613_/A vssd1 vssd1 vccd1 vccd1 _20613_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24381_ _24381_/A vssd1 vssd1 vccd1 vccd1 _27472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21593_ _21580_/X _21582_/X _21584_/X _21586_/X _21587_/X _21588_/X vssd1 vssd1 vccd1
+ vccd1 _21594_/A sky130_fd_sc_hd__mux4_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26120_ _19735_/X _26120_/D vssd1 vssd1 vccd1 vccd1 _26120_/Q sky130_fd_sc_hd__dfxtp_1
X_23332_ _23507_/A _23332_/B _23332_/C _23332_/D vssd1 vssd1 vccd1 vccd1 _23416_/B
+ sky130_fd_sc_hd__or4_1
X_20544_ _20531_/X _20533_/X _20535_/X _20537_/X _20538_/X _20539_/X vssd1 vssd1 vccd1
+ vccd1 _20545_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26051_ _26051_/CLK _26051_/D vssd1 vssd1 vccd1 vccd1 _26051_/Q sky130_fd_sc_hd__dfxtp_1
X_23263_ input51/X vssd1 vssd1 vccd1 vccd1 _23263_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20475_ _20475_/A vssd1 vssd1 vccd1 vccd1 _20475_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25002_ _25915_/Q _25981_/Q _25814_/Q _26013_/Q _24974_/X _24983_/X vssd1 vssd1 vccd1
+ vccd1 _25002_/X sky130_fd_sc_hd__mux4_1
X_22214_ _22262_/A vssd1 vssd1 vccd1 vccd1 _22214_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23194_ _23194_/A vssd1 vssd1 vccd1 vccd1 _27134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_668 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22145_ _22161_/A vssd1 vssd1 vccd1 vccd1 _22145_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22076_ _22076_/A vssd1 vssd1 vccd1 vccd1 _22076_/X sky130_fd_sc_hd__clkbuf_1
X_26953_ _22646_/X _26953_/D vssd1 vssd1 vccd1 vccd1 _26953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25904_ _27854_/CLK _25904_/D vssd1 vssd1 vccd1 vccd1 _25904_/Q sky130_fd_sc_hd__dfxtp_1
X_21027_ _21027_/A vssd1 vssd1 vccd1 vccd1 _21027_/X sky130_fd_sc_hd__clkbuf_2
X_26884_ _22400_/X _26884_/D vssd1 vssd1 vccd1 vccd1 _26884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25835_ _27850_/CLK _25835_/D vssd1 vssd1 vccd1 vccd1 _25835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13780_ _13833_/A vssd1 vssd1 vccd1 vccd1 _13780_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25766_ _17466_/X _27839_/Q _25768_/S vssd1 vssd1 vccd1 vccd1 _25767_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22978_ _25637_/A vssd1 vssd1 vccd1 vccd1 _22978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27505_ _27625_/CLK _27505_/D vssd1 vssd1 vccd1 vccd1 _27505_/Q sky130_fd_sc_hd__dfxtp_1
X_24717_ _24729_/A vssd1 vssd1 vccd1 vccd1 _24717_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21929_ _22015_/A vssd1 vssd1 vccd1 vccd1 _21997_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25697_ _25689_/X _25690_/X _25691_/X _25692_/X _25693_/X _25694_/X vssd1 vssd1 vccd1
+ vccd1 _25698_/A sky130_fd_sc_hd__mux4_1
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27436_ _27436_/CLK _27436_/D vssd1 vssd1 vccd1 vccd1 _27436_/Q sky130_fd_sc_hd__dfxtp_1
X_15450_ _15450_/A vssd1 vssd1 vccd1 vccd1 _26247_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24648_ _24648_/A vssd1 vssd1 vccd1 vccd1 _24938_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14401_ _14401_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14401_/Y sky130_fd_sc_hd__nor2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15381_ _15392_/A vssd1 vssd1 vccd1 vccd1 _15390_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27367_ _27368_/CLK _27367_/D vssd1 vssd1 vccd1 vccd1 _27367_/Q sky130_fd_sc_hd__dfxtp_1
X_24579_ _27650_/Q _24587_/B vssd1 vssd1 vccd1 vccd1 _24580_/A sky130_fd_sc_hd__and2_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _17181_/A vssd1 vssd1 vccd1 vccd1 _17120_/X sky130_fd_sc_hd__clkbuf_2
X_14332_ _26681_/Q _14322_/X _14329_/X _14331_/Y vssd1 vssd1 vccd1 vccd1 _26681_/D
+ sky130_fd_sc_hd__a31o_1
X_26318_ _20421_/X _26318_/D vssd1 vssd1 vccd1 vccd1 _26318_/Q sky130_fd_sc_hd__dfxtp_1
X_27298_ _27430_/CLK _27298_/D vssd1 vssd1 vccd1 vccd1 _27298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ input37/X vssd1 vssd1 vccd1 vccd1 _17116_/A sky130_fd_sc_hd__buf_2
X_28020__486 vssd1 vssd1 vccd1 vccd1 _28020__486/HI _28020_/A sky130_fd_sc_hd__conb_1
X_14263_ _14350_/A _14263_/B vssd1 vssd1 vccd1 vccd1 _14263_/Y sky130_fd_sc_hd__nor2_1
X_26249_ _20179_/X _26249_/D vssd1 vssd1 vccd1 vccd1 _26249_/Q sky130_fd_sc_hd__dfxtp_1
X_16002_ _16112_/A vssd1 vssd1 vccd1 vccd1 _16244_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13214_ _27339_/Q _13193_/X _13194_/X _27307_/Q _13213_/X vssd1 vssd1 vccd1 vccd1
+ _16218_/A sky130_fd_sc_hd__a221o_1
XFILLER_137_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14194_ _14220_/A vssd1 vssd1 vccd1 vccd1 _14194_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13145_ _13205_/A vssd1 vssd1 vccd1 vccd1 _13167_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_112_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17953_ _17950_/X _17952_/X _18056_/S vssd1 vssd1 vccd1 vccd1 _17953_/X sky130_fd_sc_hd__mux2_1
X_13076_ _27362_/Q _13063_/X _13064_/X _27330_/Q _13075_/X vssd1 vssd1 vccd1 vccd1
+ _13077_/A sky130_fd_sc_hd__a221o_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16904_ _16904_/A _16904_/B vssd1 vssd1 vccd1 vccd1 _16904_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_39_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater307 _27568_/CLK vssd1 vssd1 vccd1 vccd1 _27564_/CLK sky130_fd_sc_hd__clkbuf_1
X_17884_ _27795_/Q _26556_/Q _26428_/Q _26108_/Q _17782_/X _17785_/X vssd1 vssd1 vccd1
+ vccd1 _17884_/X sky130_fd_sc_hd__mux4_2
Xrepeater318 _27690_/CLK vssd1 vssd1 vccd1 vccd1 _27693_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater329 _27716_/CLK vssd1 vssd1 vccd1 vccd1 _27776_/CLK sky130_fd_sc_hd__clkbuf_1
X_19623_ _19639_/A vssd1 vssd1 vccd1 vccd1 _19623_/X sky130_fd_sc_hd__clkbuf_1
X_16835_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16835_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19554_ _26713_/Q _26681_/Q _26649_/Q _26617_/Q _18767_/X _18770_/X vssd1 vssd1 vccd1
+ vccd1 _19555_/B sky130_fd_sc_hd__mux4_2
XFILLER_202_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _14354_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16766_ _16753_/X _16763_/X _16844_/C vssd1 vssd1 vccd1 vccd1 _16766_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18505_ _26549_/Q _26517_/Q _26485_/Q _27061_/Q _17846_/X _18418_/X vssd1 vssd1 vccd1
+ vccd1 _18505_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15717_ _26131_/Q _15705_/X _15713_/X _15716_/Y vssd1 vssd1 vccd1 vccd1 _26131_/D
+ sky130_fd_sc_hd__a31o_1
X_12929_ _12929_/A _23325_/A _12929_/C _12928_/X vssd1 vssd1 vccd1 vccd1 _12933_/S
+ sky130_fd_sc_hd__or4b_4
XFILLER_94_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16697_ _16697_/A _16698_/B vssd1 vssd1 vccd1 vccd1 _16808_/A sky130_fd_sc_hd__nor2_1
X_19485_ _19485_/A vssd1 vssd1 vccd1 vccd1 _19485_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436_ _18436_/A _18322_/X vssd1 vssd1 vccd1 vccd1 _18436_/X sky130_fd_sc_hd__or2b_1
XFILLER_61_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15648_ _13116_/X _26159_/Q _15656_/S vssd1 vssd1 vccd1 vccd1 _15649_/A sky130_fd_sc_hd__mux2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15579_ _15579_/A vssd1 vssd1 vccd1 vccd1 _26190_/D sky130_fd_sc_hd__clkbuf_1
X_18367_ _18365_/X _18366_/X _18522_/S vssd1 vssd1 vccd1 vccd1 _18367_/X sky130_fd_sc_hd__mux2_2
XFILLER_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17318_ _17303_/X _17317_/X _17281_/X vssd1 vssd1 vccd1 vccd1 _17318_/X sky130_fd_sc_hd__a21bo_1
XFILLER_175_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18298_ _18455_/A vssd1 vssd1 vccd1 vccd1 _18298_/X sky130_fd_sc_hd__buf_2
XFILLER_179_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17249_ _17245_/X _17247_/X _17296_/S vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20260_ _20248_/X _20249_/X _20250_/X _20251_/X _20253_/X _20255_/X vssd1 vssd1 vccd1
+ vccd1 _20261_/A sky130_fd_sc_hd__mux4_1
XFILLER_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20191_ _20191_/A vssd1 vssd1 vccd1 vccd1 _20191_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23950_ _23997_/A vssd1 vssd1 vccd1 vccd1 _23986_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_84_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22901_ _22888_/X _22890_/X _22892_/X _22894_/X _22895_/X _22896_/X vssd1 vssd1 vccd1
+ vccd1 _22902_/A sky130_fd_sc_hd__mux4_1
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23881_ _27839_/Q _27143_/Q _25888_/Q _25856_/Q _23873_/X _23850_/X vssd1 vssd1 vccd1
+ vccd1 _23881_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25620_ _25620_/A vssd1 vssd1 vccd1 vccd1 _27789_/D sky130_fd_sc_hd__clkbuf_1
X_22832_ _22832_/A vssd1 vssd1 vccd1 vccd1 _22832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25551_ _27709_/Q _25539_/X _25540_/X vssd1 vssd1 vccd1 vccd1 _25551_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22763_ _22751_/X _22752_/X _22753_/X _22754_/X _22755_/X _22756_/X vssd1 vssd1 vccd1
+ vccd1 _22764_/A sky130_fd_sc_hd__mux4_1
XFILLER_198_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24502_ _24403_/A _24633_/C _24501_/X _24499_/X vssd1 vssd1 vccd1 vccd1 _27521_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ _21714_/A vssd1 vssd1 vccd1 vccd1 _21714_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25482_ _25456_/X _25461_/X _25462_/X _24859_/B _25463_/X vssd1 vssd1 vccd1 vccd1
+ _25482_/X sky130_fd_sc_hd__o311a_1
X_22694_ _22694_/A vssd1 vssd1 vccd1 vccd1 _22694_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27221_ _27222_/CLK _27221_/D vssd1 vssd1 vccd1 vccd1 _27221_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24433_ _27616_/Q _24433_/B vssd1 vssd1 vccd1 vccd1 _24434_/A sky130_fd_sc_hd__and2_1
X_21645_ _21631_/X _21632_/X _21633_/X _21634_/X _21635_/X _21636_/X vssd1 vssd1 vccd1
+ vccd1 _21646_/A sky130_fd_sc_hd__mux4_1
XFILLER_200_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27152_ _27153_/CLK _27152_/D vssd1 vssd1 vccd1 vccd1 _27152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24364_ _27564_/Q _24372_/B vssd1 vssd1 vccd1 vccd1 _24365_/A sky130_fd_sc_hd__and2_1
XANTENNA_50 _18061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21576_ _21576_/A vssd1 vssd1 vccd1 vccd1 _21576_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_61 _18289_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _18451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26103_ _19675_/X _26103_/D vssd1 vssd1 vccd1 vccd1 _26103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23315_ input70/X vssd1 vssd1 vccd1 vccd1 _23315_/Y sky130_fd_sc_hd__inv_2
X_27083_ _27083_/CLK _27083_/D vssd1 vssd1 vccd1 vccd1 _27083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_83 _18850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20527_ _20527_/A vssd1 vssd1 vccd1 vccd1 _20527_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_94 _19180_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24295_ _16274_/X _16276_/Y _16277_/Y _24279_/A vssd1 vssd1 vccd1 vccd1 _27426_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_181_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26034_ _27850_/CLK _26034_/D vssd1 vssd1 vccd1 vccd1 _26034_/Q sky130_fd_sc_hd__dfxtp_1
X_23246_ _17514_/X _27158_/Q _23248_/S vssd1 vssd1 vccd1 vccd1 _23247_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20458_ _20445_/X _20447_/X _20449_/X _20451_/X _20452_/X _20453_/X vssd1 vssd1 vccd1
+ vccd1 _20459_/A sky130_fd_sc_hd__mux4_1
XFILLER_106_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23177_ _23177_/A vssd1 vssd1 vccd1 vccd1 _27127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20389_ _20389_/A vssd1 vssd1 vccd1 vccd1 _20389_/X sky130_fd_sc_hd__clkbuf_1
X_22128_ _22176_/A vssd1 vssd1 vccd1 vccd1 _22128_/X sky130_fd_sc_hd__clkbuf_1
X_27985_ _27985_/A _15897_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
XFILLER_88_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14950_ _14950_/A vssd1 vssd1 vccd1 vccd1 _26461_/D sky130_fd_sc_hd__clkbuf_1
X_22059_ _22051_/X _22052_/X _22053_/X _22054_/X _22055_/X _22056_/X vssd1 vssd1 vccd1
+ vccd1 _22060_/A sky130_fd_sc_hd__mux4_1
X_26936_ _22586_/X _26936_/D vssd1 vssd1 vccd1 vccd1 _26936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13901_ _26826_/Q _13893_/X _13899_/X _13900_/Y vssd1 vssd1 vccd1 vccd1 _26826_/D
+ sky130_fd_sc_hd__a31o_1
X_14881_ _26491_/Q _13417_/X _14883_/S vssd1 vssd1 vccd1 vccd1 _14882_/A sky130_fd_sc_hd__mux2_1
X_26867_ _22342_/X _26867_/D vssd1 vssd1 vccd1 vccd1 _26867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13832_ _13844_/A vssd1 vssd1 vccd1 vccd1 _13832_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16620_ _16660_/A _16618_/B _16619_/X vssd1 vssd1 vccd1 vccd1 _16620_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25818_ _26017_/CLK _25818_/D vssd1 vssd1 vccd1 vccd1 _25818_/Q sky130_fd_sc_hd__dfxtp_1
X_26798_ _22098_/X _26798_/D vssd1 vssd1 vccd1 vccd1 _26798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16551_ _16826_/A _16552_/B vssd1 vssd1 vccd1 vccd1 _16551_/Y sky130_fd_sc_hd__nor2_1
X_13763_ _13779_/A vssd1 vssd1 vccd1 vccd1 _13847_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25749_ _17440_/X _27831_/Q _25757_/S vssd1 vssd1 vccd1 vccd1 _25750_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15502_ _15502_/A vssd1 vssd1 vccd1 vccd1 _26224_/D sky130_fd_sc_hd__clkbuf_1
X_19270_ _19428_/A vssd1 vssd1 vccd1 vccd1 _19409_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_71_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16482_ _16482_/A _16482_/B _16481_/X vssd1 vssd1 vccd1 vccd1 _16483_/A sky130_fd_sc_hd__or3b_1
X_13694_ _26900_/Q _13682_/X _13692_/X _13693_/Y vssd1 vssd1 vccd1 vccd1 _26900_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18221_ _26953_/Q _26921_/Q _26889_/Q _26857_/Q _17999_/X _18000_/X vssd1 vssd1 vccd1
+ vccd1 _18221_/X sky130_fd_sc_hd__mux4_2
X_15433_ _15433_/A vssd1 vssd1 vccd1 vccd1 _26255_/D sky130_fd_sc_hd__clkbuf_1
X_27419_ _27675_/CLK _27419_/D vssd1 vssd1 vccd1 vccd1 _27419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18152_ _26950_/Q _26918_/Q _26886_/Q _26854_/Q _18101_/X _18129_/X vssd1 vssd1 vccd1
+ vccd1 _18152_/X sky130_fd_sc_hd__mux4_2
XFILLER_15_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15364_ _14750_/X _26285_/Q _15368_/S vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14315_ _26687_/Q _14310_/X _14311_/X _14314_/Y vssd1 vssd1 vccd1 vccd1 _26687_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17103_ _27202_/Q _17102_/X _17128_/S vssd1 vssd1 vccd1 vccd1 _17104_/A sky130_fd_sc_hd__mux2_1
X_18083_ _26691_/Q _26659_/Q _26627_/Q _26595_/Q _18004_/X _18005_/X vssd1 vssd1 vccd1
+ vccd1 _18084_/A sky130_fd_sc_hd__mux4_2
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15295_ _26315_/Q _13366_/X _15295_/S vssd1 vssd1 vccd1 vccd1 _15296_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17034_ _16998_/X _17032_/X _17033_/X vssd1 vssd1 vccd1 vccd1 _17034_/X sky130_fd_sc_hd__a21bo_1
X_14246_ _14333_/A _14248_/B vssd1 vssd1 vccd1 vccd1 _14246_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14177_ _14354_/A _14187_/B vssd1 vssd1 vccd1 vccd1 _14177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _14750_/A vssd1 vssd1 vccd1 vccd1 _13128_/X sky130_fd_sc_hd__buf_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _26527_/Q _26495_/Q _26463_/Q _27039_/Q _18984_/X _18863_/X vssd1 vssd1 vccd1
+ vccd1 _18985_/X sky130_fd_sc_hd__mux4_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17936_ _17936_/A _17935_/X vssd1 vssd1 vccd1 vccd1 _17936_/X sky130_fd_sc_hd__or2b_1
X_13059_ _27064_/Q _13058_/X _13079_/S vssd1 vssd1 vccd1 vccd1 _13060_/A sky130_fd_sc_hd__mux2_1
Xrepeater104 _25901_/CLK vssd1 vssd1 vccd1 vccd1 _27155_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater115 _27686_/CLK vssd1 vssd1 vccd1 vccd1 _27299_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater126 _26038_/CLK vssd1 vssd1 vccd1 vccd1 _26037_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater137 _27095_/CLK vssd1 vssd1 vccd1 vccd1 _27094_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17867_ _17867_/A _17813_/X vssd1 vssd1 vccd1 vccd1 _17867_/X sky130_fd_sc_hd__or2b_1
Xrepeater148 _27420_/CLK vssd1 vssd1 vccd1 vccd1 _26040_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater159 _27407_/CLK vssd1 vssd1 vccd1 vccd1 _25878_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19606_ _19638_/A vssd1 vssd1 vccd1 vccd1 _19606_/X sky130_fd_sc_hd__clkbuf_1
X_16818_ _16697_/A _16499_/A _16809_/Y _16809_/A _16817_/Y vssd1 vssd1 vccd1 vccd1
+ _16818_/X sky130_fd_sc_hd__a32o_1
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17798_ _18474_/A vssd1 vssd1 vccd1 vccd1 _18322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19537_ _26968_/Q _26936_/Q _26904_/Q _26872_/Q _18824_/X _18826_/X vssd1 vssd1 vccd1
+ vccd1 _19537_/X sky130_fd_sc_hd__mux4_1
X_16749_ _16751_/A _16749_/B vssd1 vssd1 vccd1 vccd1 _16765_/D sky130_fd_sc_hd__xnor2_1
XFILLER_185_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ _19466_/X _19467_/X _19468_/S vssd1 vssd1 vccd1 vccd1 _19468_/X sky130_fd_sc_hd__mux2_2
XFILLER_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18419_ _26545_/Q _26513_/Q _26481_/Q _27057_/Q _18392_/X _18418_/X vssd1 vssd1 vccd1
+ vccd1 _18419_/X sky130_fd_sc_hd__mux4_1
XFILLER_195_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19399_ _19399_/A vssd1 vssd1 vccd1 vccd1 _19399_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21430_ _21478_/A vssd1 vssd1 vccd1 vccd1 _21430_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21361_ _21377_/A vssd1 vssd1 vccd1 vccd1 _21361_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23100_ _23100_/A vssd1 vssd1 vccd1 vccd1 _27093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20312_ _20302_/X _20303_/X _20304_/X _20305_/X _20306_/X _20307_/X vssd1 vssd1 vccd1
+ vccd1 _20313_/A sky130_fd_sc_hd__mux4_1
Xinput70 la1_oenb[7] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_6
XFILLER_135_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24080_ _27389_/Q _24084_/B vssd1 vssd1 vccd1 vccd1 _24081_/A sky130_fd_sc_hd__and2_1
X_21292_ _21292_/A vssd1 vssd1 vccd1 vccd1 _21292_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23031_ _23025_/X _23026_/X _23027_/X _23028_/X _23029_/X _23030_/X vssd1 vssd1 vccd1
+ vccd1 _23032_/A sky130_fd_sc_hd__mux4_1
X_20243_ _20243_/A vssd1 vssd1 vccd1 vccd1 _20243_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20174_ _20162_/X _20163_/X _20164_/X _20165_/X _20167_/X _20169_/X vssd1 vssd1 vccd1
+ vccd1 _20175_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27770_ _27770_/CLK _27770_/D vssd1 vssd1 vccd1 vccd1 _27770_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24982_ _27827_/Q _27131_/Q _25876_/Q _25844_/Q _24972_/X _23638_/B vssd1 vssd1 vccd1
+ vccd1 _24982_/X sky130_fd_sc_hd__mux4_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26721_ _21836_/X _26721_/D vssd1 vssd1 vccd1 vccd1 _26721_/Q sky130_fd_sc_hd__dfxtp_1
X_23933_ _23931_/X _23932_/X _23940_/S vssd1 vssd1 vccd1 vccd1 _23933_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26652_ _21594_/X _26652_/D vssd1 vssd1 vccd1 vccd1 _26652_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23864_ _23864_/A vssd1 vssd1 vccd1 vccd1 _23864_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25603_ _25572_/X _25582_/X _25583_/X _24962_/B _25584_/X vssd1 vssd1 vccd1 vccd1
+ _25603_/X sky130_fd_sc_hd__o311a_1
X_22815_ _22802_/X _22804_/X _22806_/X _22808_/X _22809_/X _22810_/X vssd1 vssd1 vccd1
+ vccd1 _22816_/A sky130_fd_sc_hd__mux4_1
XFILLER_199_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26583_ _21354_/X _26583_/D vssd1 vssd1 vccd1 vccd1 _26583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23795_ _23793_/X _23794_/X _23795_/S vssd1 vssd1 vccd1 vccd1 _23795_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25534_ _25564_/A vssd1 vssd1 vccd1 vccd1 _25534_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22746_ _22746_/A vssd1 vssd1 vccd1 vccd1 _22746_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25465_ _25438_/X _25151_/B _25464_/X _25452_/X vssd1 vssd1 vccd1 vccd1 _25465_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_160_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22677_ _22665_/X _22666_/X _22667_/X _22668_/X _22669_/X _22670_/X vssd1 vssd1 vccd1
+ vccd1 _22678_/A sky130_fd_sc_hd__mux4_1
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27204_ _27353_/CLK _27204_/D vssd1 vssd1 vccd1 vccd1 _27204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24416_ _27588_/Q _24422_/B vssd1 vssd1 vccd1 vccd1 _24417_/A sky130_fd_sc_hd__and2_1
X_21628_ _21628_/A vssd1 vssd1 vccd1 vccd1 _21628_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25396_ _27737_/Q input48/X _25402_/S vssd1 vssd1 vccd1 vccd1 _25397_/A sky130_fd_sc_hd__mux2_1
X_27135_ _27135_/CLK _27135_/D vssd1 vssd1 vccd1 vccd1 _27135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24347_ _24347_/A vssd1 vssd1 vccd1 vccd1 _27456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21559_ _21545_/X _21546_/X _21547_/X _21548_/X _21549_/X _21550_/X vssd1 vssd1 vccd1
+ vccd1 _21560_/A sky130_fd_sc_hd__mux4_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14100_ _14127_/A vssd1 vssd1 vccd1 vccd1 _14112_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15080_ _15080_/A vssd1 vssd1 vccd1 vccd1 _26411_/D sky130_fd_sc_hd__clkbuf_1
X_27066_ _27408_/CLK _27066_/D vssd1 vssd1 vccd1 vccd1 _27066_/Q sky130_fd_sc_hd__dfxtp_1
X_24278_ _16202_/X _16204_/Y _16206_/X _24273_/X vssd1 vssd1 vccd1 vccd1 _27415_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_101_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_868 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14031_ _14503_/A vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26017_ _26017_/CLK _26017_/D vssd1 vssd1 vccd1 vccd1 _26017_/Q sky130_fd_sc_hd__dfxtp_1
X_23229_ _17488_/X _27150_/Q _23237_/S vssd1 vssd1 vccd1 vccd1 _23230_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18770_ _19486_/A vssd1 vssd1 vccd1 vccd1 _18770_/X sky130_fd_sc_hd__clkbuf_2
X_15982_ _15985_/A vssd1 vssd1 vccd1 vccd1 _15982_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27968_ _27968_/A _15867_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17721_ _27422_/Q vssd1 vssd1 vccd1 vccd1 _17721_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26919_ _22518_/X _26919_/D vssd1 vssd1 vccd1 vccd1 _26919_/Q sky130_fd_sc_hd__dfxtp_1
X_14933_ _14933_/A vssd1 vssd1 vccd1 vccd1 _26469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17652_ _17495_/X _25897_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _17653_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14864_ _26499_/Q _13392_/X _14868_/S vssd1 vssd1 vccd1 vccd1 _14865_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _16603_/A _16793_/A vssd1 vssd1 vccd1 vccd1 _16604_/B sky130_fd_sc_hd__xnor2_1
X_13815_ _13908_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13815_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17583_ _17583_/A vssd1 vssd1 vccd1 vccd1 _25866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14795_ _16224_/A vssd1 vssd1 vccd1 vccd1 _14795_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19322_ _27813_/Q _26574_/Q _26446_/Q _26126_/Q _19255_/X _19321_/X vssd1 vssd1 vccd1
+ vccd1 _19322_/X sky130_fd_sc_hd__mux4_2
X_13746_ _13926_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13746_/Y sky130_fd_sc_hd__nor2_1
X_16534_ _16534_/A _16534_/B vssd1 vssd1 vccd1 vccd1 _16535_/B sky130_fd_sc_hd__xor2_1
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19253_ _19412_/A vssd1 vssd1 vccd1 vccd1 _19253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13677_ _13691_/A vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16465_ _16392_/Y _16399_/Y _16433_/Y _16464_/X vssd1 vssd1 vccd1 vccd1 _16482_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ _18198_/X _18200_/X _18202_/X _18203_/X vssd1 vssd1 vccd1 vccd1 _18204_/X
+ sky130_fd_sc_hd__o211a_1
X_15416_ _26262_/Q _13331_/X _15418_/S vssd1 vssd1 vccd1 vccd1 _15417_/A sky130_fd_sc_hd__mux2_1
X_19184_ _27807_/Q _26568_/Q _26440_/Q _26120_/Q _19118_/X _19183_/X vssd1 vssd1 vccd1
+ vccd1 _19184_/X sky130_fd_sc_hd__mux4_2
X_16396_ _16745_/B _16396_/B vssd1 vssd1 vccd1 vccd1 _16396_/X sky130_fd_sc_hd__and2_1
XFILLER_185_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18135_ _18057_/X _18132_/X _18134_/X _18062_/X vssd1 vssd1 vccd1 vccd1 _18135_/X
+ sky130_fd_sc_hd__o211a_1
X_15347_ _15347_/A vssd1 vssd1 vccd1 vccd1 _26293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_781 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15278_ _26323_/Q _13341_/X _15284_/S vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__mux2_1
X_18066_ _18322_/A vssd1 vssd1 vccd1 vccd1 _18066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14229_ _26717_/Q _14225_/X _14220_/X _14228_/Y vssd1 vssd1 vccd1 vccd1 _26717_/D
+ sky130_fd_sc_hd__a31o_1
X_17017_ input35/X vssd1 vssd1 vccd1 vccd1 _17266_/A sky130_fd_sc_hd__buf_2
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18968_ _26815_/Q _26783_/Q _26751_/Q _26719_/Q _18870_/X _18967_/X vssd1 vssd1 vccd1
+ vccd1 _18969_/B sky130_fd_sc_hd__mux4_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _17919_/A vssd1 vssd1 vccd1 vccd1 _25946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18899_ _26941_/Q _26909_/Q _26877_/Q _26845_/Q _18896_/X _18898_/X vssd1 vssd1 vccd1
+ vccd1 _18899_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20930_ _20930_/A vssd1 vssd1 vccd1 vccd1 _20930_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20861_ _20861_/A vssd1 vssd1 vccd1 vccd1 _20861_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22600_ _22600_/A vssd1 vssd1 vccd1 vccd1 _22600_/X sky130_fd_sc_hd__clkbuf_1
X_23580_ _23600_/A vssd1 vssd1 vccd1 vccd1 _23595_/S sky130_fd_sc_hd__clkbuf_2
X_20792_ _20792_/A vssd1 vssd1 vccd1 vccd1 _22540_/A sky130_fd_sc_hd__buf_4
XFILLER_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22531_ _22519_/X _22520_/X _22521_/X _22522_/X _22524_/X _22526_/X vssd1 vssd1 vccd1
+ vccd1 _22532_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25250_ _25250_/A _25241_/A vssd1 vssd1 vccd1 vccd1 _25250_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22462_ _22462_/A vssd1 vssd1 vccd1 vccd1 _22462_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24201_ _24201_/A vssd1 vssd1 vccd1 vccd1 _27369_/D sky130_fd_sc_hd__clkbuf_1
X_21413_ _21585_/A vssd1 vssd1 vccd1 vccd1 _21478_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25181_ _25181_/A _25181_/B vssd1 vssd1 vccd1 vccd1 _25182_/B sky130_fd_sc_hd__xnor2_1
X_22393_ _22385_/X _22386_/X _22387_/X _22388_/X _22389_/X _22390_/X vssd1 vssd1 vccd1
+ vccd1 _22394_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24132_ _27444_/Q _24140_/B vssd1 vssd1 vccd1 vccd1 _24133_/A sky130_fd_sc_hd__and2_1
X_21344_ _21392_/A vssd1 vssd1 vccd1 vccd1 _21344_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24063_ _24063_/A vssd1 vssd1 vccd1 vccd1 _24072_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21275_ _21269_/X _21270_/X _21271_/X _21272_/X _21273_/X _21274_/X vssd1 vssd1 vccd1
+ vccd1 _21276_/A sky130_fd_sc_hd__mux4_1
X_23014_ _23030_/A vssd1 vssd1 vccd1 vccd1 _23014_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20226_ _20216_/X _20217_/X _20218_/X _20219_/X _20220_/X _20221_/X vssd1 vssd1 vccd1
+ vccd1 _20227_/A sky130_fd_sc_hd__mux4_1
XFILLER_103_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27822_ _25728_/X _27822_/D vssd1 vssd1 vccd1 vccd1 _27822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20157_ _20157_/A vssd1 vssd1 vccd1 vccd1 _20157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27753_ _27753_/CLK _27753_/D vssd1 vssd1 vccd1 vccd1 _27753_/Q sky130_fd_sc_hd__dfxtp_1
X_24965_ _24965_/A _24965_/B vssd1 vssd1 vccd1 vccd1 _24966_/B sky130_fd_sc_hd__or2_1
XFILLER_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ _20076_/X _20077_/X _20078_/X _20079_/X _20081_/X _20083_/X vssd1 vssd1 vccd1
+ vccd1 _20089_/A sky130_fd_sc_hd__mux4_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26704_ _21776_/X _26704_/D vssd1 vssd1 vccd1 vccd1 _26704_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23916_ _27082_/Q _27114_/Q _23939_/S vssd1 vssd1 vccd1 vccd1 _23916_/X sky130_fd_sc_hd__mux2_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27684_ _27684_/CLK _27684_/D vssd1 vssd1 vccd1 vccd1 _27975_/A sky130_fd_sc_hd__dfxtp_1
X_24896_ _27769_/Q _27768_/Q _24896_/C vssd1 vssd1 vccd1 vccd1 _24902_/B sky130_fd_sc_hd__and3_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26635_ _21536_/X _26635_/D vssd1 vssd1 vccd1 vccd1 _26635_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23847_ _27075_/Q _23812_/X _23813_/X _27107_/Q _23814_/X vssd1 vssd1 vccd1 vccd1
+ _23847_/X sky130_fd_sc_hd__a221o_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13870_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13600_/Y sky130_fd_sc_hd__nor2_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _15741_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14580_/Y sky130_fd_sc_hd__nor2_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26566_ _21294_/X _26566_/D vssd1 vssd1 vccd1 vccd1 _26566_/Q sky130_fd_sc_hd__dfxtp_1
X_23778_ _27828_/Q _27132_/Q _25877_/Q _25845_/Q _23777_/X _23744_/X vssd1 vssd1 vccd1
+ vccd1 _23778_/X sky130_fd_sc_hd__mux4_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _27346_/Q _13529_/X _13530_/X _27314_/Q _13169_/X vssd1 vssd1 vccd1 vccd1
+ _14493_/A sky130_fd_sc_hd__a221oi_4
XFILLER_14_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25517_ _25517_/A vssd1 vssd1 vccd1 vccd1 _25517_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22729_ _22716_/X _22718_/X _22720_/X _22722_/X _22723_/X _22724_/X vssd1 vssd1 vccd1
+ vccd1 _22730_/A sky130_fd_sc_hd__mux4_1
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26497_ _21052_/X _26497_/D vssd1 vssd1 vccd1 vccd1 _26497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _27390_/Q _16132_/A _16137_/X _26056_/Q _16249_/X vssd1 vssd1 vccd1 vccd1
+ _24287_/A sky130_fd_sc_hd__a221o_1
XFILLER_201_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _15773_/A vssd1 vssd1 vccd1 vccd1 _13792_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_25448_ _25539_/A vssd1 vssd1 vccd1 vccd1 _25448_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15201_ _14724_/X _26357_/Q _15201_/S vssd1 vssd1 vccd1 vccd1 _15202_/A sky130_fd_sc_hd__mux2_1
X_16181_ _16201_/A vssd1 vssd1 vccd1 vccd1 _16215_/B sky130_fd_sc_hd__clkbuf_1
X_25379_ _25379_/A vssd1 vssd1 vccd1 vccd1 _27729_/D sky130_fd_sc_hd__clkbuf_1
X_13393_ _26979_/Q _13392_/X _13399_/S vssd1 vssd1 vccd1 vccd1 _13394_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _26388_/Q _13337_/X _15140_/S vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__mux2_1
X_27118_ _27299_/CLK _27118_/D vssd1 vssd1 vccd1 vccd1 _27118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19940_ _19988_/A vssd1 vssd1 vccd1 vccd1 _19940_/X sky130_fd_sc_hd__clkbuf_1
X_15063_ _15063_/A vssd1 vssd1 vccd1 vccd1 _26419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27049_ _22972_/X _27049_/D vssd1 vssd1 vccd1 vccd1 _27049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14014_ _14381_/A _14029_/B vssd1 vssd1 vccd1 vccd1 _14014_/Y sky130_fd_sc_hd__nor2_1
X_19871_ _19887_/A vssd1 vssd1 vccd1 vccd1 _19871_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18822_ _18814_/X _18819_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _18822_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18753_ _26037_/Q _17763_/X _18757_/S vssd1 vssd1 vccd1 vccd1 _18754_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15965_ _15967_/A vssd1 vssd1 vccd1 vccd1 _15965_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17704_ _17704_/A vssd1 vssd1 vccd1 vccd1 _25920_/D sky130_fd_sc_hd__clkbuf_1
X_14916_ _14753_/X _26476_/Q _14918_/S vssd1 vssd1 vccd1 vccd1 _14917_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18684_ _18684_/A vssd1 vssd1 vccd1 vccd1 _26006_/D sky130_fd_sc_hd__clkbuf_1
X_15896_ _15899_/A vssd1 vssd1 vccd1 vccd1 _15896_/Y sky130_fd_sc_hd__inv_2
X_17635_ _17635_/A vssd1 vssd1 vccd1 vccd1 _25889_/D sky130_fd_sc_hd__clkbuf_1
X_14847_ _14847_/A vssd1 vssd1 vccd1 vccd1 _26507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17566_ _17566_/A vssd1 vssd1 vccd1 vccd1 _25858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14778_ _14778_/A vssd1 vssd1 vccd1 vccd1 _26533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19305_ _26285_/Q _26253_/Q _26221_/Q _26189_/Q _19297_/X _18930_/A vssd1 vssd1 vccd1
+ vccd1 _19305_/X sky130_fd_sc_hd__mux4_2
X_16517_ _16805_/B vssd1 vssd1 vccd1 vccd1 _16824_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13729_ _26887_/Q _13724_/X _13718_/X _13728_/Y vssd1 vssd1 vccd1 vccd1 _26887_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17497_ _17497_/A vssd1 vssd1 vccd1 vccd1 _25833_/D sky130_fd_sc_hd__clkbuf_1
X_19236_ _26154_/Q _26090_/Q _27018_/Q _26986_/Q _19165_/X _19188_/X vssd1 vssd1 vccd1
+ vccd1 _19237_/B sky130_fd_sc_hd__mux4_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16448_ _16446_/Y _16447_/Y _25910_/Q vssd1 vssd1 vccd1 vccd1 _16449_/B sky130_fd_sc_hd__a21oi_1
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19167_ _19261_/A _19167_/B vssd1 vssd1 vccd1 vccd1 _19167_/X sky130_fd_sc_hd__or2_1
XFILLER_192_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16379_ _16388_/A _16447_/B _16357_/A _16744_/A _16360_/A vssd1 vssd1 vccd1 vccd1
+ _16380_/B sky130_fd_sc_hd__o41a_1
XFILLER_185_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18118_ _26532_/Q _26500_/Q _26468_/Q _27044_/Q _18117_/X _17986_/X vssd1 vssd1 vccd1
+ vccd1 _18118_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19098_ _26276_/Q _26244_/Q _26212_/Q _26180_/Q _19028_/X _19074_/X vssd1 vssd1 vccd1
+ vccd1 _19098_/X sky130_fd_sc_hd__mux4_2
XFILLER_172_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18049_ _26401_/Q _26369_/Q _26337_/Q _26305_/Q _18048_/X _17943_/X vssd1 vssd1 vccd1
+ vccd1 _18049_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21060_ _21126_/A vssd1 vssd1 vccd1 vccd1 _21060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20011_ _20077_/A vssd1 vssd1 vccd1 vccd1 _20011_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24750_ _24750_/A _24759_/B vssd1 vssd1 vccd1 vccd1 _24750_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21962_ _21962_/A vssd1 vssd1 vccd1 vccd1 _21962_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23701_ _24925_/A _27255_/Q _23705_/S vssd1 vssd1 vccd1 vccd1 _23702_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20913_ _20905_/X _20906_/X _20907_/X _20908_/X _20909_/X _20910_/X vssd1 vssd1 vccd1
+ vccd1 _20914_/A sky130_fd_sc_hd__mux4_1
X_24681_ _27174_/Q _24685_/B vssd1 vssd1 vccd1 vccd1 _24681_/X sky130_fd_sc_hd__or2_1
X_21893_ _21879_/X _21880_/X _21881_/X _21882_/X _21883_/X _21884_/X vssd1 vssd1 vccd1
+ vccd1 _21894_/A sky130_fd_sc_hd__mux4_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23632_ _25102_/S vssd1 vssd1 vccd1 vccd1 _25004_/S sky130_fd_sc_hd__buf_2
X_26420_ _20779_/X _26420_/D vssd1 vssd1 vccd1 vccd1 _26420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20844_ _20832_/X _20833_/X _20834_/X _20835_/X _20836_/X _20837_/X vssd1 vssd1 vccd1
+ vccd1 _20845_/A sky130_fd_sc_hd__mux4_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26351_ _20543_/X _26351_/D vssd1 vssd1 vccd1 vccd1 _26351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23563_ _23600_/A vssd1 vssd1 vccd1 vccd1 _23576_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20775_ _20852_/A vssd1 vssd1 vccd1 vccd1 _20775_/X sky130_fd_sc_hd__clkbuf_2
X_25302_ _25310_/A _27511_/Q vssd1 vssd1 vccd1 vccd1 _25304_/A sky130_fd_sc_hd__or2_1
X_22514_ _22514_/A vssd1 vssd1 vccd1 vccd1 _22514_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26282_ _20297_/X _26282_/D vssd1 vssd1 vccd1 vccd1 _26282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23494_ input29/X _23482_/X _23493_/X _23487_/X vssd1 vssd1 vccd1 vccd1 _27190_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28021_ _28021_/A _15982_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
X_25233_ _27535_/Q _27503_/Q vssd1 vssd1 vccd1 vccd1 _25250_/A sky130_fd_sc_hd__and2_1
XFILLER_7_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22445_ _22433_/X _22434_/X _22435_/X _22436_/X _22438_/X _22440_/X vssd1 vssd1 vccd1
+ vccd1 _22446_/A sky130_fd_sc_hd__mux4_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25164_ _25164_/A _25164_/B vssd1 vssd1 vccd1 vccd1 _25165_/B sky130_fd_sc_hd__nor2_1
X_22376_ _22376_/A vssd1 vssd1 vccd1 vccd1 _22376_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24115_ _27405_/Q _24117_/B vssd1 vssd1 vccd1 vccd1 _24116_/A sky130_fd_sc_hd__and2_1
XFILLER_159_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21327_ _21585_/A vssd1 vssd1 vccd1 vccd1 _21392_/A sky130_fd_sc_hd__clkbuf_2
X_25095_ _27080_/Q _27112_/Q _25102_/S vssd1 vssd1 vccd1 vccd1 _25095_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24046_ _27097_/Q _27129_/Q _24046_/S vssd1 vssd1 vccd1 vccd1 _24046_/X sky130_fd_sc_hd__mux2_1
X_21258_ _21290_/A vssd1 vssd1 vccd1 vccd1 _21258_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_563 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20209_ _20209_/A vssd1 vssd1 vccd1 vccd1 _20209_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21189_ _21179_/X _21180_/X _21181_/X _21182_/X _21183_/X _21184_/X vssd1 vssd1 vccd1
+ vccd1 _21190_/A sky130_fd_sc_hd__mux4_1
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27805_ _25670_/X _27805_/D vssd1 vssd1 vccd1 vccd1 _27805_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25997_ _27122_/CLK _25997_/D vssd1 vssd1 vccd1 vccd1 _25997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _26119_/Q _15747_/X _15740_/X _15749_/Y vssd1 vssd1 vccd1 vccd1 _26119_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _12962_/A vssd1 vssd1 vccd1 vccd1 _27816_/D sky130_fd_sc_hd__clkbuf_1
X_27736_ _27748_/CLK _27736_/D vssd1 vssd1 vccd1 vccd1 _27736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24948_ _24954_/C _24948_/B vssd1 vssd1 vccd1 vccd1 _24949_/B sky130_fd_sc_hd__or2_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _15775_/A _14707_/B vssd1 vssd1 vccd1 vccd1 _14701_/Y sky130_fd_sc_hd__nor2_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_310 _18080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27667_ _27667_/CLK _27667_/D vssd1 vssd1 vccd1 vccd1 _27667_/Q sky130_fd_sc_hd__dfxtp_1
X_15681_ _13204_/X _26144_/Q _15689_/S vssd1 vssd1 vccd1 vccd1 _15682_/A sky130_fd_sc_hd__mux2_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24879_ _27652_/Q _24861_/X _24878_/Y _24864_/X vssd1 vssd1 vccd1 vccd1 _27652_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _19062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _23035_/A _17420_/B _23033_/A _23035_/C vssd1 vssd1 vccd1 vccd1 _24003_/A
+ sky130_fd_sc_hd__and4_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_332 _25733_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26618_ _21472_/X _26618_/D vssd1 vssd1 vccd1 vccd1 _26618_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _26583_/Q _14630_/X _14624_/X _14631_/Y vssd1 vssd1 vccd1 vccd1 _26583_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_343 _13350_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_354 _14531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_365 _26813_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27598_ _27601_/CLK _27598_/D vssd1 vssd1 vccd1 vccd1 _27598_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _17338_/X _17351_/B vssd1 vssd1 vccd1 vccd1 _17351_/X sky130_fd_sc_hd__and2b_1
X_14563_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14563_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26549_ _21228_/X _26549_/D vssd1 vssd1 vccd1 vccd1 _26549_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16833_/A _16576_/B vssd1 vssd1 vccd1 vccd1 _16595_/B sky130_fd_sc_hd__nor2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _26953_/Q _13510_/X _13505_/X _13513_/Y vssd1 vssd1 vccd1 vccd1 _26953_/D
+ sky130_fd_sc_hd__a31o_1
X_14494_ _15754_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _14494_/Y sky130_fd_sc_hd__nor2_1
X_17282_ _17242_/X _17280_/X _17281_/X vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__a21bo_1
XFILLER_202_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19021_ _19018_/X _19020_/X _19047_/S vssd1 vssd1 vccd1 vccd1 _19021_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ _16134_/A vssd1 vssd1 vccd1 vccd1 _13868_/A sky130_fd_sc_hd__clkbuf_2
X_16233_ _26051_/Q _16233_/B _16233_/C vssd1 vssd1 vccd1 vccd1 _16233_/X sky130_fd_sc_hd__and3_1
XFILLER_201_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13376_ _14766_/A vssd1 vssd1 vccd1 vccd1 _13376_/X sky130_fd_sc_hd__clkbuf_4
X_16164_ _27530_/Q _16242_/S vssd1 vssd1 vccd1 vccd1 _16164_/X sky130_fd_sc_hd__or2b_1
XFILLER_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15115_ _15115_/A vssd1 vssd1 vccd1 vccd1 _26395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16095_ _16313_/B _16313_/C _16457_/B vssd1 vssd1 vccd1 vccd1 _16310_/A sky130_fd_sc_hd__a21oi_1
XFILLER_141_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19923_ _20270_/A vssd1 vssd1 vccd1 vccd1 _19990_/A sky130_fd_sc_hd__clkbuf_2
X_15046_ _15335_/A _15262_/B vssd1 vssd1 vccd1 vccd1 _15103_/A sky130_fd_sc_hd__or2_4
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19854_ _19886_/A vssd1 vssd1 vccd1 vccd1 _19854_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18805_ _19299_/A vssd1 vssd1 vccd1 vccd1 _19555_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19785_ _19801_/A vssd1 vssd1 vccd1 vccd1 _19785_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16997_ input36/X vssd1 vssd1 vccd1 vccd1 _17303_/A sky130_fd_sc_hd__buf_2
X_18736_ _18736_/A vssd1 vssd1 vccd1 vccd1 _26029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _15949_/A vssd1 vssd1 vccd1 vccd1 _15948_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18667_ _18667_/A vssd1 vssd1 vccd1 vccd1 _25998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ _15881_/A vssd1 vssd1 vccd1 vccd1 _15879_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _17618_/A vssd1 vssd1 vccd1 vccd1 _25881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18598_ _18613_/A _18598_/B vssd1 vssd1 vccd1 vccd1 _25113_/A sky130_fd_sc_hd__nand2_1
X_17549_ _17450_/X _25851_/Q _17551_/S vssd1 vssd1 vccd1 vccd1 _17550_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20560_ _20550_/X _20551_/X _20552_/X _20553_/X _20554_/X _20555_/X vssd1 vssd1 vccd1
+ vccd1 _20561_/A sky130_fd_sc_hd__mux4_1
XFILLER_165_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19219_ _18814_/X _19218_/X _18785_/X vssd1 vssd1 vccd1 vccd1 _19219_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20491_ _20491_/A vssd1 vssd1 vccd1 vccd1 _20491_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22230_ _22262_/A vssd1 vssd1 vccd1 vccd1 _22230_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22161_ _22161_/A vssd1 vssd1 vccd1 vccd1 _22161_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21112_ _21128_/A vssd1 vssd1 vccd1 vccd1 _21112_/X sky130_fd_sc_hd__clkbuf_1
X_22092_ _22092_/A vssd1 vssd1 vccd1 vccd1 _22092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25920_ _25986_/CLK _25920_/D vssd1 vssd1 vccd1 vccd1 _25920_/Q sky130_fd_sc_hd__dfxtp_1
X_21043_ _21215_/A vssd1 vssd1 vccd1 vccd1 _21113_/A sky130_fd_sc_hd__buf_2
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25851_ _25884_/CLK _25851_/D vssd1 vssd1 vccd1 vccd1 _25851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24802_ _27633_/Q _24798_/X _24800_/Y _24801_/X vssd1 vssd1 vccd1 vccd1 _27633_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25782_ _17488_/X _27846_/Q _25790_/S vssd1 vssd1 vccd1 vccd1 _25783_/A sky130_fd_sc_hd__mux2_1
X_22994_ _25636_/A vssd1 vssd1 vccd1 vccd1 _22994_/X sky130_fd_sc_hd__clkbuf_1
X_27521_ _27523_/CLK _27521_/D vssd1 vssd1 vccd1 vccd1 _27521_/Q sky130_fd_sc_hd__dfxtp_1
X_21945_ _21930_/X _21932_/X _21934_/X _21936_/X _21937_/X _21938_/X vssd1 vssd1 vccd1
+ vccd1 _21946_/A sky130_fd_sc_hd__mux4_1
XFILLER_27_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24733_ _24733_/A _24748_/A vssd1 vssd1 vccd1 vccd1 _24733_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24664_ _24635_/A _24660_/X _24662_/X _24663_/X vssd1 vssd1 vccd1 vccd1 _27583_/D
+ sky130_fd_sc_hd__o211a_1
X_27452_ _27452_/CLK _27452_/D vssd1 vssd1 vccd1 vccd1 _27452_/Q sky130_fd_sc_hd__dfxtp_1
X_21876_ _21876_/A vssd1 vssd1 vccd1 vccd1 _21876_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26403_ _20719_/X _26403_/D vssd1 vssd1 vccd1 vccd1 _26403_/Q sky130_fd_sc_hd__dfxtp_1
X_23615_ _27782_/Q vssd1 vssd1 vccd1 vccd1 _24960_/A sky130_fd_sc_hd__buf_2
XFILLER_199_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20827_ _20827_/A vssd1 vssd1 vccd1 vccd1 _20827_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24595_ _24595_/A vssd1 vssd1 vccd1 vccd1 _27557_/D sky130_fd_sc_hd__clkbuf_1
X_27383_ _27383_/CLK _27383_/D vssd1 vssd1 vccd1 vccd1 _27383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26334_ _20479_/X _26334_/D vssd1 vssd1 vccd1 vccd1 _26334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23546_ _23623_/S vssd1 vssd1 vccd1 vccd1 _23559_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20758_ _20758_/A vssd1 vssd1 vccd1 vccd1 _20758_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26265_ _20239_/X _26265_/D vssd1 vssd1 vccd1 vccd1 _26265_/Q sky130_fd_sc_hd__dfxtp_1
X_23477_ input22/X _23469_/X _23476_/X _23474_/X vssd1 vssd1 vccd1 vccd1 _27183_/D
+ sky130_fd_sc_hd__o211a_1
X_20689_ _20758_/A vssd1 vssd1 vccd1 vccd1 _20689_/X sky130_fd_sc_hd__clkbuf_2
X_28004_ _28004_/A _15875_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
X_25216_ _27533_/Q _27501_/Q vssd1 vssd1 vccd1 vccd1 _25218_/A sky130_fd_sc_hd__nand2_1
X_13230_ _13230_/A vssd1 vssd1 vccd1 vccd1 _27036_/D sky130_fd_sc_hd__clkbuf_1
X_22428_ _22428_/A vssd1 vssd1 vccd1 vccd1 _22428_/X sky130_fd_sc_hd__clkbuf_1
X_26196_ _20001_/X _26196_/D vssd1 vssd1 vccd1 vccd1 _26196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_614 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13161_ _14769_/A vssd1 vssd1 vccd1 vccd1 _13161_/X sky130_fd_sc_hd__buf_2
X_25147_ _25147_/A _25146_/X vssd1 vssd1 vccd1 vccd1 _25150_/A sky130_fd_sc_hd__or2b_1
X_22359_ _22347_/X _22348_/X _22349_/X _22350_/X _22352_/X _22354_/X vssd1 vssd1 vccd1
+ vccd1 _22360_/A sky130_fd_sc_hd__mux4_1
XFILLER_152_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25078_ _27838_/Q _27142_/Q _25887_/Q _25855_/Q _25061_/X _24975_/X vssd1 vssd1 vccd1
+ vccd1 _25078_/X sky130_fd_sc_hd__mux4_1
XFILLER_123_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13092_ _27296_/Q _13142_/B vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__and2_2
XFILLER_152_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24029_ _27855_/Q _27159_/Q _25904_/Q _25872_/Q _24014_/X _23991_/X vssd1 vssd1 vccd1
+ vccd1 _24029_/X sky130_fd_sc_hd__mux4_1
X_16920_ _24264_/A _24263_/A _24255_/A _24261_/A vssd1 vssd1 vccd1 vccd1 _25583_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16851_ _16851_/A _16851_/B vssd1 vssd1 vccd1 vccd1 _16852_/B sky130_fd_sc_hd__or2_1
XFILLER_120_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15802_ _15802_/A vssd1 vssd1 vccd1 vccd1 _26098_/D sky130_fd_sc_hd__clkbuf_1
X_19570_ _19637_/A vssd1 vssd1 vccd1 vccd1 _19570_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16782_ _16778_/Y _16781_/X _16768_/X vssd1 vssd1 vccd1 vccd1 _16782_/X sky130_fd_sc_hd__a21o_1
X_13994_ _16277_/A vssd1 vssd1 vccd1 vccd1 _14367_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18521_ _26422_/Q _26390_/Q _26358_/Q _26326_/Q _17959_/A _17904_/X vssd1 vssd1 vccd1
+ vccd1 _18521_/X sky130_fd_sc_hd__mux4_1
X_15733_ _26125_/Q _15721_/X _15727_/X _15732_/Y vssd1 vssd1 vccd1 vccd1 _26125_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27719_ _27719_/CLK _27719_/D vssd1 vssd1 vccd1 vccd1 _27719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12945_/A vssd1 vssd1 vccd1 vccd1 _27823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18452_ _26835_/Q _26803_/Q _26771_/Q _26739_/Q _18085_/X _17913_/X vssd1 vssd1 vccd1
+ vccd1 _18452_/X sky130_fd_sc_hd__mux4_2
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _15664_/A vssd1 vssd1 vccd1 vccd1 _26152_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _25106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _13190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17403_ input3/X vssd1 vssd1 vccd1 vccd1 _25641_/A sky130_fd_sc_hd__buf_6
XANTENNA_173 _16298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ _14671_/A vssd1 vssd1 vccd1 vccd1 _14615_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _16277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18383_ _18383_/A _18317_/X vssd1 vssd1 vccd1 vccd1 _18383_/X sky130_fd_sc_hd__or2b_1
XFILLER_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _26182_/Q _16240_/A _15595_/S vssd1 vssd1 vccd1 vccd1 _15596_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _16442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17332_/X _17333_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17334_/X sky130_fd_sc_hd__mux2_2
XFILLER_53_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14546_ _15708_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17265_ _27847_/Q _27151_/Q _25896_/Q _25864_/Q _17264_/X _17252_/X vssd1 vssd1 vccd1
+ vccd1 _17265_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14477_ _26634_/Q _14460_/X _14474_/X _14476_/Y vssd1 vssd1 vccd1 vccd1 _26634_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19004_ _19004_/A _19004_/B vssd1 vssd1 vccd1 vccd1 _19004_/X sky130_fd_sc_hd__or2_1
X_16216_ _27380_/Q vssd1 vssd1 vccd1 vccd1 _17674_/B sky130_fd_sc_hd__clkinv_2
X_13428_ _13456_/A vssd1 vssd1 vccd1 vccd1 _13583_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17196_ _17181_/X _17195_/X _17159_/X vssd1 vssd1 vccd1 vccd1 _17196_/X sky130_fd_sc_hd__a21bo_1
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16147_ _16797_/A vssd1 vssd1 vccd1 vccd1 _16798_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13359_ _13359_/A vssd1 vssd1 vccd1 vccd1 _26990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16078_ _16593_/A vssd1 vssd1 vccd1 vccd1 _16648_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15029_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15029_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19906_ _19898_/X _19899_/X _19900_/X _19901_/X _19903_/X _19905_/X vssd1 vssd1 vccd1
+ vccd1 _19907_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19837_ _19901_/A vssd1 vssd1 vccd1 vccd1 _19837_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19768_ _19800_/A vssd1 vssd1 vccd1 vccd1 _19768_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18719_ _18719_/A vssd1 vssd1 vccd1 vccd1 _26021_/D sky130_fd_sc_hd__clkbuf_1
X_19699_ _19715_/A vssd1 vssd1 vccd1 vccd1 _19699_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21730_ _21730_/A vssd1 vssd1 vccd1 vccd1 _21730_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21661_ _21647_/X _21648_/X _21649_/X _21650_/X _21652_/X _21654_/X vssd1 vssd1 vccd1
+ vccd1 _21662_/A sky130_fd_sc_hd__mux4_1
XFILLER_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23400_ _27762_/Q vssd1 vssd1 vccd1 vccd1 _24756_/A sky130_fd_sc_hd__inv_2
X_20612_ _20598_/X _20599_/X _20600_/X _20601_/X _20603_/X _20605_/X vssd1 vssd1 vccd1
+ vccd1 _20613_/A sky130_fd_sc_hd__mux4_1
XFILLER_178_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24380_ _27577_/Q _24380_/B vssd1 vssd1 vccd1 vccd1 _24381_/A sky130_fd_sc_hd__and2_1
XFILLER_71_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21592_ _21592_/A vssd1 vssd1 vccd1 vccd1 _21592_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_812 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23331_ _23331_/A _23331_/B _23331_/C _23331_/D vssd1 vssd1 vccd1 vccd1 _23332_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20543_ _20543_/A vssd1 vssd1 vccd1 vccd1 _20543_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26050_ _26051_/CLK _26050_/D vssd1 vssd1 vccd1 vccd1 _26050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23262_ _27747_/Q vssd1 vssd1 vccd1 vccd1 _23262_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20474_ _20464_/X _20465_/X _20466_/X _20467_/X _20468_/X _20469_/X vssd1 vssd1 vccd1
+ vccd1 _20475_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25001_ _27829_/Q _27133_/Q _25878_/Q _25846_/Q _24972_/X _24991_/X vssd1 vssd1 vccd1
+ vccd1 _25001_/X sky130_fd_sc_hd__mux4_1
X_22213_ _22261_/A vssd1 vssd1 vccd1 vccd1 _22213_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23193_ _17437_/X _27134_/Q _23193_/S vssd1 vssd1 vccd1 vccd1 _23194_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_422 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22144_ _22176_/A vssd1 vssd1 vccd1 vccd1 _22144_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22075_ _22067_/X _22068_/X _22069_/X _22070_/X _22071_/X _22072_/X vssd1 vssd1 vccd1
+ vccd1 _22076_/A sky130_fd_sc_hd__mux4_1
X_26952_ _22644_/X _26952_/D vssd1 vssd1 vccd1 vccd1 _26952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25903_ _27155_/CLK _25903_/D vssd1 vssd1 vccd1 vccd1 _25903_/Q sky130_fd_sc_hd__dfxtp_1
X_21026_ _21042_/A vssd1 vssd1 vccd1 vccd1 _21026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26883_ _22398_/X _26883_/D vssd1 vssd1 vccd1 vccd1 _26883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25834_ _26001_/CLK _25834_/D vssd1 vssd1 vccd1 vccd1 _25834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25765_ _25765_/A vssd1 vssd1 vccd1 vccd1 _27838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22977_ _25657_/A vssd1 vssd1 vccd1 vccd1 _25637_/A sky130_fd_sc_hd__clkbuf_2
X_27504_ _27625_/CLK _27504_/D vssd1 vssd1 vccd1 vccd1 _27504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24716_ _27187_/Q _24725_/B vssd1 vssd1 vccd1 vccd1 _24716_/X sky130_fd_sc_hd__or2_1
X_21928_ _21928_/A vssd1 vssd1 vccd1 vccd1 _21928_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25696_ _25696_/A vssd1 vssd1 vccd1 vccd1 _25696_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27435_ _27435_/CLK _27435_/D vssd1 vssd1 vccd1 vccd1 _27435_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21859_ _21844_/X _21846_/X _21848_/X _21850_/X _21851_/X _21852_/X vssd1 vssd1 vccd1
+ vccd1 _21860_/A sky130_fd_sc_hd__mux4_1
XFILLER_188_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24647_ _24828_/A _24828_/B vssd1 vssd1 vccd1 vccd1 _24648_/A sky130_fd_sc_hd__and2_1
XFILLER_163_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14400_ _26656_/Q _14392_/X _14398_/X _14399_/Y vssd1 vssd1 vccd1 vccd1 _26656_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15380_/A vssd1 vssd1 vccd1 vccd1 _26278_/D sky130_fd_sc_hd__clkbuf_1
X_27366_ _27443_/CLK _27366_/D vssd1 vssd1 vccd1 vccd1 _27366_/Q sky130_fd_sc_hd__dfxtp_2
X_24578_ _24589_/A vssd1 vssd1 vccd1 vccd1 _24587_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_156_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14331_ _14331_/A _14335_/B vssd1 vssd1 vccd1 vccd1 _14331_/Y sky130_fd_sc_hd__nor2_1
X_26317_ _20419_/X _26317_/D vssd1 vssd1 vccd1 vccd1 _26317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23529_ _23623_/S vssd1 vssd1 vccd1 vccd1 _23542_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27297_ _27425_/CLK _27297_/D vssd1 vssd1 vccd1 vccd1 _27297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ _26707_/Q _14256_/X _14258_/X _14261_/Y vssd1 vssd1 vccd1 vccd1 _26707_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_167_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17050_ _17050_/A vssd1 vssd1 vccd1 vccd1 _27919_/A sky130_fd_sc_hd__clkbuf_1
X_26248_ _20177_/X _26248_/D vssd1 vssd1 vccd1 vccd1 _26248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16001_ _16001_/A _16001_/B _16001_/C _16001_/D vssd1 vssd1 vccd1 vccd1 _16112_/A
+ sky130_fd_sc_hd__and4_1
X_13213_ _27275_/Q _13237_/B vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__and2_1
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ _26731_/Q _14186_/X _14181_/X _14192_/Y vssd1 vssd1 vccd1 vccd1 _26731_/D
+ sky130_fd_sc_hd__a31o_1
X_26179_ _19939_/X _26179_/D vssd1 vssd1 vccd1 vccd1 _26179_/Q sky130_fd_sc_hd__dfxtp_1
X_13144_ _14759_/A vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__buf_2
XFILLER_48_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17952_ _26942_/Q _26910_/Q _26878_/Q _26846_/Q _17922_/X _17951_/X vssd1 vssd1 vccd1
+ vccd1 _17952_/X sky130_fd_sc_hd__mux4_2
X_13075_ _27298_/Q _13109_/B vssd1 vssd1 vccd1 vccd1 _13075_/X sky130_fd_sc_hd__and2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16903_ _16879_/A _16879_/B _16878_/B _16599_/Y vssd1 vssd1 vccd1 vccd1 _16904_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater308 _27468_/CLK vssd1 vssd1 vccd1 vccd1 _27568_/CLK sky130_fd_sc_hd__clkbuf_1
X_17883_ _24611_/A vssd1 vssd1 vccd1 vccd1 _18028_/A sky130_fd_sc_hd__clkbuf_1
Xrepeater319 _27760_/CLK vssd1 vssd1 vccd1 vccd1 _27766_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19622_ _19638_/A vssd1 vssd1 vccd1 vccd1 _19622_/X sky130_fd_sc_hd__clkbuf_1
X_16834_ _16800_/C _16832_/X _16833_/Y vssd1 vssd1 vccd1 vccd1 _16834_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19553_ _19551_/X _19552_/X _19553_/S vssd1 vssd1 vccd1 vccd1 _19553_/X sky130_fd_sc_hd__mux2_1
X_16765_ _16765_/A _16765_/B _16765_/C _16765_/D vssd1 vssd1 vccd1 vccd1 _16844_/C
+ sky130_fd_sc_hd__or4_1
X_13977_ _14032_/A vssd1 vssd1 vccd1 vccd1 _13992_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18504_ _18437_/X _18503_/X _18483_/X vssd1 vssd1 vccd1 vccd1 _18504_/X sky130_fd_sc_hd__o21a_1
X_15716_ _15716_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15716_/Y sky130_fd_sc_hd__nor2_1
X_12928_ _12928_/A _12928_/B _12928_/C _12928_/D vssd1 vssd1 vccd1 vccd1 _12928_/X
+ sky130_fd_sc_hd__and4_1
X_19484_ _19524_/A _19484_/B vssd1 vssd1 vccd1 vccd1 _19484_/X sky130_fd_sc_hd__or2_1
X_16696_ _27392_/Q _16094_/X _16412_/X _25960_/Q _16495_/Y vssd1 vssd1 vccd1 vccd1
+ _16698_/B sky130_fd_sc_hd__a221o_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18435_ _26162_/Q _26098_/Q _27026_/Q _26994_/Q _18298_/X _18387_/X vssd1 vssd1 vccd1
+ vccd1 _18436_/A sky130_fd_sc_hd__mux4_2
XFILLER_34_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15647_ _15693_/S vssd1 vssd1 vccd1 vccd1 _15656_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18366_ _26415_/Q _26383_/Q _26351_/Q _26319_/Q _17903_/X _17904_/X vssd1 vssd1 vccd1
+ vccd1 _18366_/X sky130_fd_sc_hd__mux4_1
X_15578_ _26190_/Q _14747_/A _15584_/S vssd1 vssd1 vccd1 vccd1 _15579_/A sky130_fd_sc_hd__mux2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17317_ _25836_/Q _26035_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__mux2_1
X_14529_ _26619_/Q _14514_/X _14426_/B _14528_/Y vssd1 vssd1 vccd1 vccd1 _26619_/D
+ sky130_fd_sc_hd__a31o_1
X_18297_ _17995_/X _18291_/X _18293_/X _18295_/X _18352_/S vssd1 vssd1 vccd1 vccd1
+ _18309_/B sky130_fd_sc_hd__a221o_1
XFILLER_30_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17248_ input38/X vssd1 vssd1 vccd1 vccd1 _17296_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17179_ _25926_/Q _25992_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17180_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20190_ _20181_/X _20183_/X _20185_/X _20187_/X _20188_/X _20189_/X vssd1 vssd1 vccd1
+ vccd1 _20191_/A sky130_fd_sc_hd__mux4_1
XFILLER_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22900_ _22900_/A vssd1 vssd1 vccd1 vccd1 _22900_/X sky130_fd_sc_hd__clkbuf_1
X_23880_ _23849_/X _23878_/X _23879_/X _23864_/X vssd1 vssd1 vccd1 vccd1 _27283_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22831_ _22821_/X _22822_/X _22823_/X _22824_/X _22825_/X _22826_/X vssd1 vssd1 vccd1
+ vccd1 _22832_/A sky130_fd_sc_hd__mux4_1
XFILLER_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25550_ _24782_/A _25534_/X _25546_/Y _25549_/X _25527_/X vssd1 vssd1 vccd1 vccd1
+ _27772_/D sky130_fd_sc_hd__a221oi_1
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22762_ _22762_/A vssd1 vssd1 vccd1 vccd1 _22762_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21713_ _21705_/X _21706_/X _21707_/X _21708_/X _21709_/X _21710_/X vssd1 vssd1 vccd1
+ vccd1 _21714_/A sky130_fd_sc_hd__mux4_1
X_24501_ _27587_/Q _24505_/B vssd1 vssd1 vccd1 vccd1 _24501_/X sky130_fd_sc_hd__or2_1
X_25481_ _27697_/Q _25479_/X _25480_/X vssd1 vssd1 vccd1 vccd1 _25481_/Y sky130_fd_sc_hd__a21oi_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22693_ _22681_/X _22682_/X _22683_/X _22684_/X _22685_/X _22686_/X vssd1 vssd1 vccd1
+ vccd1 _22694_/A sky130_fd_sc_hd__mux4_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27220_ _27224_/CLK _27220_/D vssd1 vssd1 vccd1 vccd1 _27220_/Q sky130_fd_sc_hd__dfxtp_1
X_21644_ _21644_/A vssd1 vssd1 vccd1 vccd1 _21644_/X sky130_fd_sc_hd__clkbuf_1
X_24432_ _24432_/A vssd1 vssd1 vccd1 vccd1 _27494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27151_ _27151_/CLK _27151_/D vssd1 vssd1 vccd1 vccd1 _27151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24363_ _24363_/A vssd1 vssd1 vccd1 vccd1 _24372_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_178_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21575_ _21561_/X _21562_/X _21563_/X _21564_/X _21566_/X _21568_/X vssd1 vssd1 vccd1
+ vccd1 _21576_/A sky130_fd_sc_hd__mux4_1
XANTENNA_40 _18000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_51 _18084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_62 _18293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23314_ _27730_/Q _23305_/Y _23255_/Y input48/X _23313_/X vssd1 vssd1 vccd1 vccd1
+ _23320_/B sky130_fd_sc_hd__o221ai_1
X_26102_ _19673_/X _26102_/D vssd1 vssd1 vccd1 vccd1 _26102_/Q sky130_fd_sc_hd__dfxtp_1
X_27082_ _27115_/CLK _27082_/D vssd1 vssd1 vccd1 vccd1 _27082_/Q sky130_fd_sc_hd__dfxtp_1
X_20526_ _20512_/X _20513_/X _20514_/X _20515_/X _20517_/X _20519_/X vssd1 vssd1 vccd1
+ vccd1 _20527_/A sky130_fd_sc_hd__mux4_1
XANTENNA_73 _18480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24294_ _16268_/X _16270_/Y _16271_/X _24279_/X vssd1 vssd1 vccd1 vccd1 _27425_/D
+ sky130_fd_sc_hd__o31a_1
XANTENNA_84 _18868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_95 _19209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23245_ _23245_/A vssd1 vssd1 vccd1 vccd1 _27157_/D sky130_fd_sc_hd__clkbuf_1
X_26033_ _27151_/CLK _26033_/D vssd1 vssd1 vccd1 vccd1 _26033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20457_ _20457_/A vssd1 vssd1 vccd1 vccd1 _20457_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23176_ _27127_/Q _17769_/X _23176_/S vssd1 vssd1 vccd1 vccd1 _23177_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20388_ _20376_/X _20377_/X _20378_/X _20379_/X _20380_/X _20381_/X vssd1 vssd1 vccd1
+ vccd1 _20389_/A sky130_fd_sc_hd__mux4_1
XFILLER_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22127_ _22175_/A vssd1 vssd1 vccd1 vccd1 _22127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_414 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27984_ _27984_/A _15898_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
XFILLER_133_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22058_ _22058_/A vssd1 vssd1 vccd1 vccd1 _22058_/X sky130_fd_sc_hd__clkbuf_1
X_26935_ _22584_/X _26935_/D vssd1 vssd1 vccd1 vccd1 _26935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13900_ _13900_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21009_ _21041_/A vssd1 vssd1 vccd1 vccd1 _21009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26866_ _22340_/X _26866_/D vssd1 vssd1 vccd1 vccd1 _26866_/Q sky130_fd_sc_hd__dfxtp_1
X_14880_ _14880_/A vssd1 vssd1 vccd1 vccd1 _26492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13831_ _26849_/Q _13819_/X _13820_/X _13830_/Y vssd1 vssd1 vccd1 vccd1 _26849_/D
+ sky130_fd_sc_hd__a31o_1
X_25817_ _27414_/CLK _25817_/D vssd1 vssd1 vccd1 vccd1 _25817_/Q sky130_fd_sc_hd__dfxtp_1
X_26797_ _22096_/X _26797_/D vssd1 vssd1 vccd1 vccd1 _26797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16550_ _16824_/B _16550_/B vssd1 vssd1 vccd1 vccd1 _16550_/X sky130_fd_sc_hd__and2b_1
X_13762_ _15695_/D _13762_/B vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__or2_2
X_25748_ _25805_/S vssd1 vssd1 vccd1 vccd1 _25757_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _13111_/X _26224_/Q _15501_/S vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16481_ _16481_/A _16464_/X vssd1 vssd1 vccd1 vccd1 _16481_/X sky130_fd_sc_hd__or2b_1
X_13693_ _13874_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13693_/Y sky130_fd_sc_hd__nor2_1
X_25679_ _25673_/X _25674_/X _25675_/X _25676_/X _25677_/X _25678_/X vssd1 vssd1 vccd1
+ vccd1 _25680_/A sky130_fd_sc_hd__mux4_1
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18220_ _27808_/Q _26569_/Q _26441_/Q _26121_/Q _17996_/X _17997_/X vssd1 vssd1 vccd1
+ vccd1 _18220_/X sky130_fd_sc_hd__mux4_2
X_27418_ _27418_/CLK _27418_/D vssd1 vssd1 vccd1 vccd1 _27418_/Q sky130_fd_sc_hd__dfxtp_1
X_15432_ _26255_/Q _13353_/X _15440_/S vssd1 vssd1 vccd1 vccd1 _15433_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18151_ _27805_/Q _26566_/Q _26438_/Q _26118_/Q _18099_/X _18126_/X vssd1 vssd1 vccd1
+ vccd1 _18151_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15363_ _15363_/A vssd1 vssd1 vccd1 vccd1 _26286_/D sky130_fd_sc_hd__clkbuf_1
X_27349_ _27350_/CLK _27349_/D vssd1 vssd1 vccd1 vccd1 _27349_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17102_ _17100_/X _17101_/X _17113_/S vssd1 vssd1 vccd1 vccd1 _17102_/X sky130_fd_sc_hd__mux2_1
X_14314_ _14401_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14314_/Y sky130_fd_sc_hd__nor2_1
X_18082_ _18079_/X _18080_/X _18514_/S vssd1 vssd1 vccd1 vccd1 _18082_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15294_ _15294_/A vssd1 vssd1 vccd1 vccd1 _26316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033_ _17220_/A vssd1 vssd1 vccd1 vccd1 _17033_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14245_ _26713_/Q _14238_/X _14242_/X _14244_/Y vssd1 vssd1 vccd1 vccd1 _26713_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14176_ _14215_/A vssd1 vssd1 vccd1 vccd1 _14187_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13127_ _13127_/A vssd1 vssd1 vccd1 vccd1 _14750_/A sky130_fd_sc_hd__clkbuf_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _19414_/A vssd1 vssd1 vccd1 vccd1 _18984_/X sky130_fd_sc_hd__buf_2
XFILLER_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _18322_/A vssd1 vssd1 vccd1 vccd1 _17935_/X sky130_fd_sc_hd__clkbuf_1
X_13058_ _14715_/A vssd1 vssd1 vccd1 vccd1 _13058_/X sky130_fd_sc_hd__buf_2
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater105 _25900_/CLK vssd1 vssd1 vccd1 vccd1 _25901_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater116 _27285_/CLK vssd1 vssd1 vccd1 vccd1 _27686_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater127 _25941_/CLK vssd1 vssd1 vccd1 vccd1 _26007_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater138 _26026_/CLK vssd1 vssd1 vccd1 vccd1 _27842_/CLK sky130_fd_sc_hd__clkbuf_1
X_17866_ _26683_/Q _26651_/Q _26619_/Q _26587_/Q _17865_/X _17810_/X vssd1 vssd1 vccd1
+ vccd1 _17867_/A sky130_fd_sc_hd__mux4_1
XFILLER_61_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater149 _27420_/CLK vssd1 vssd1 vccd1 vccd1 _27857_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16817_ _14756_/A _16501_/X _16098_/X _25961_/Q _16490_/Y vssd1 vssd1 vccd1 vccd1
+ _16817_/Y sky130_fd_sc_hd__a221oi_2
X_19605_ _19637_/A vssd1 vssd1 vccd1 vccd1 _19605_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17797_ _27595_/Q vssd1 vssd1 vccd1 vccd1 _18474_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19536_ _19431_/X _19535_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _19536_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_548 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16748_ _16744_/Y _16746_/X _16765_/A vssd1 vssd1 vccd1 vccd1 _16748_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19467_ _26548_/Q _26516_/Q _26484_/Q _27060_/Q _19401_/X _19445_/X vssd1 vssd1 vccd1
+ vccd1 _19467_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16679_ _16715_/C _16393_/Y _16738_/B _16877_/A vssd1 vssd1 vccd1 vccd1 _16679_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_62_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18418_ _18418_/A vssd1 vssd1 vccd1 vccd1 _18418_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19398_ _19351_/X _19397_/X _19354_/X vssd1 vssd1 vccd1 vccd1 _19398_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _26414_/Q _26382_/Q _26350_/Q _26318_/Q _18085_/A _18141_/A vssd1 vssd1 vccd1
+ vccd1 _18349_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21360_ _21392_/A vssd1 vssd1 vccd1 vccd1 _21360_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20311_ _20311_/A vssd1 vssd1 vccd1 vccd1 _20311_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput60 la1_oenb[27] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_6
X_21291_ _21285_/X _21286_/X _21287_/X _21288_/X _21289_/X _21290_/X vssd1 vssd1 vccd1
+ vccd1 _21292_/A sky130_fd_sc_hd__mux4_1
Xinput71 la1_oenb[8] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_2
X_23030_ _23030_/A vssd1 vssd1 vccd1 vccd1 _23030_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20242_ _20232_/X _20233_/X _20234_/X _20235_/X _20236_/X _20237_/X vssd1 vssd1 vccd1
+ vccd1 _20243_/A sky130_fd_sc_hd__mux4_1
XFILLER_104_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20173_ _20173_/A vssd1 vssd1 vccd1 vccd1 _20173_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24981_ _24981_/A vssd1 vssd1 vccd1 vccd1 _27672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26720_ _21834_/X _26720_/D vssd1 vssd1 vccd1 vccd1 _26720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23932_ _27084_/Q _27116_/Q _23939_/S vssd1 vssd1 vccd1 vccd1 _23932_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26651_ _21592_/X _26651_/D vssd1 vssd1 vccd1 vccd1 _26651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23863_ _27076_/Q _23860_/X _23861_/X _27108_/Q _23862_/X vssd1 vssd1 vccd1 vccd1
+ _23863_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25602_ _25599_/X _25600_/Y _25601_/Y _25446_/X vssd1 vssd1 vccd1 vccd1 _27781_/D
+ sky130_fd_sc_hd__a211oi_1
X_22814_ _22814_/A vssd1 vssd1 vccd1 vccd1 _22814_/X sky130_fd_sc_hd__clkbuf_1
X_26582_ _21352_/X _26582_/D vssd1 vssd1 vccd1 vccd1 _26582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23794_ _25916_/Q _25982_/Q _25815_/Q _26014_/Q _23747_/X _23786_/X vssd1 vssd1 vccd1
+ vccd1 _23794_/X sky130_fd_sc_hd__mux4_1
XFILLER_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25533_ _24776_/A _25504_/X _25529_/Y _25532_/X _25527_/X vssd1 vssd1 vccd1 vccd1
+ _27769_/D sky130_fd_sc_hd__a221oi_1
X_22745_ _22735_/X _22736_/X _22737_/X _22738_/X _22739_/X _22740_/X vssd1 vssd1 vccd1
+ vccd1 _22746_/A sky130_fd_sc_hd__mux4_1
XFILLER_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22676_ _22676_/A vssd1 vssd1 vccd1 vccd1 _22676_/X sky130_fd_sc_hd__clkbuf_1
X_25464_ _25456_/X _25461_/X _25462_/X _24846_/B _25463_/X vssd1 vssd1 vccd1 vccd1
+ _25464_/X sky130_fd_sc_hd__o311a_1
XFILLER_185_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27203_ _27350_/CLK _27203_/D vssd1 vssd1 vccd1 vccd1 _27203_/Q sky130_fd_sc_hd__dfxtp_1
X_21627_ _21615_/X _21616_/X _21617_/X _21618_/X _21619_/X _21620_/X vssd1 vssd1 vccd1
+ vccd1 _21628_/A sky130_fd_sc_hd__mux4_1
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24415_ _24415_/A vssd1 vssd1 vccd1 vccd1 _27486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25395_ _25395_/A vssd1 vssd1 vccd1 vccd1 _27736_/D sky130_fd_sc_hd__clkbuf_1
X_27134_ _27412_/CLK _27134_/D vssd1 vssd1 vccd1 vccd1 _27134_/Q sky130_fd_sc_hd__dfxtp_1
X_21558_ _21558_/A vssd1 vssd1 vccd1 vccd1 _21558_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24346_ _27556_/Q _24350_/B vssd1 vssd1 vccd1 vccd1 _24347_/A sky130_fd_sc_hd__and2_1
XFILLER_181_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20509_ _20509_/A vssd1 vssd1 vccd1 vccd1 _20509_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24277_ _16209_/X _16211_/Y _16212_/X _24273_/X vssd1 vssd1 vccd1 vccd1 _27414_/D
+ sky130_fd_sc_hd__o31a_1
X_27065_ _23032_/X _27065_/D vssd1 vssd1 vccd1 vccd1 _27065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21489_ _21475_/X _21476_/X _21477_/X _21478_/X _21480_/X _21482_/X vssd1 vssd1 vccd1
+ vccd1 _21490_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14030_ _26787_/Q _14024_/X _14019_/X _14029_/Y vssd1 vssd1 vccd1 vccd1 _26787_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_10_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23228_ _23239_/A vssd1 vssd1 vccd1 vccd1 _23237_/S sky130_fd_sc_hd__buf_2
XFILLER_153_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26016_ _26016_/CLK _26016_/D vssd1 vssd1 vccd1 vccd1 _26016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23159_ _27119_/Q _17744_/X _23165_/S vssd1 vssd1 vccd1 vccd1 _23160_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15981_ _15985_/A vssd1 vssd1 vccd1 vccd1 _15981_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27967_ _27967_/A _15866_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ _17720_/A vssd1 vssd1 vccd1 vccd1 _25925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26918_ _22516_/X _26918_/D vssd1 vssd1 vccd1 vccd1 _26918_/Q sky130_fd_sc_hd__dfxtp_1
X_14932_ _14775_/X _26469_/Q _14940_/S vssd1 vssd1 vccd1 vccd1 _14933_/A sky130_fd_sc_hd__mux2_1
X_17651_ _17651_/A vssd1 vssd1 vccd1 vccd1 _25896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26849_ _22278_/X _26849_/D vssd1 vssd1 vccd1 vccd1 _26849_/Q sky130_fd_sc_hd__dfxtp_1
X_14863_ _14863_/A vssd1 vssd1 vccd1 vccd1 _26500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16602_ _16602_/A _16602_/B vssd1 vssd1 vccd1 vccd1 _16793_/A sky130_fd_sc_hd__or2_1
X_13814_ _13827_/A vssd1 vssd1 vccd1 vccd1 _13825_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_1163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17582_ _17498_/X _25866_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17583_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ _14794_/A vssd1 vssd1 vccd1 vccd1 _26528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19321_ _19321_/A vssd1 vssd1 vccd1 vccd1 _19321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16533_ _16292_/B _16292_/C _16802_/A _16106_/A vssd1 vssd1 vccd1 vccd1 _16534_/B
+ sky130_fd_sc_hd__o31a_1
X_13745_ _13745_/A vssd1 vssd1 vccd1 vccd1 _13745_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19252_ _19158_/X _19251_/X _19229_/X vssd1 vssd1 vccd1 vccd1 _19252_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16464_ _16686_/A _16450_/Y _16610_/A _16692_/C vssd1 vssd1 vccd1 vccd1 _16464_/X
+ sky130_fd_sc_hd__and4bb_1
X_13676_ _13759_/B vssd1 vssd1 vccd1 vccd1 _13676_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18203_ _18384_/A vssd1 vssd1 vccd1 vccd1 _18203_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15415_ _15415_/A vssd1 vssd1 vccd1 vccd1 _26263_/D sky130_fd_sc_hd__clkbuf_1
X_19183_ _19321_/A vssd1 vssd1 vccd1 vccd1 _19183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16395_ _16395_/A _16395_/B vssd1 vssd1 vccd1 vccd1 _16395_/Y sky130_fd_sc_hd__nand2_1
X_18134_ _18134_/A _17978_/X vssd1 vssd1 vccd1 vccd1 _18134_/X sky130_fd_sc_hd__or2b_1
XFILLER_106_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15346_ _14724_/X _26293_/Q _15346_/S vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_793 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18065_ _26146_/Q _26082_/Q _27010_/Q _26978_/Q _18041_/X _17959_/X vssd1 vssd1 vccd1
+ vccd1 _18067_/A sky130_fd_sc_hd__mux4_1
X_15277_ _15277_/A vssd1 vssd1 vccd1 vccd1 _26324_/D sky130_fd_sc_hd__clkbuf_1
X_17016_ _27827_/Q _27131_/Q _25876_/Q _25844_/Q _17015_/X _16989_/X vssd1 vssd1 vccd1
+ vccd1 _17016_/X sky130_fd_sc_hd__mux4_1
X_14228_ _14406_/A _14234_/B vssd1 vssd1 vccd1 vccd1 _14228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _26743_/Q _14157_/X _14151_/X _14158_/Y vssd1 vssd1 vccd1 vccd1 _26743_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _19486_/A vssd1 vssd1 vccd1 vccd1 _18967_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _18028_/A _17918_/B _17918_/C vssd1 vssd1 vccd1 vccd1 _17919_/A sky130_fd_sc_hd__and3_1
X_18898_ _19445_/A vssd1 vssd1 vccd1 vccd1 _18898_/X sky130_fd_sc_hd__buf_4
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17849_ _26394_/Q _26362_/Q _26330_/Q _26298_/Q _17846_/X _17848_/X vssd1 vssd1 vccd1
+ vccd1 _17849_/X sky130_fd_sc_hd__mux4_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20860_ _20848_/X _20849_/X _20850_/X _20851_/X _20852_/X _20853_/X vssd1 vssd1 vccd1
+ vccd1 _20861_/A sky130_fd_sc_hd__mux4_1
XFILLER_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ _26967_/Q _26935_/Q _26903_/Q _26871_/Q _18824_/X _19412_/X vssd1 vssd1 vccd1
+ vccd1 _19519_/X sky130_fd_sc_hd__mux4_1
XFILLER_179_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20791_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20791_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22530_ _22530_/A vssd1 vssd1 vccd1 vccd1 _22530_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22461_ _22452_/X _22454_/X _22456_/X _22458_/X _22459_/X _22460_/X vssd1 vssd1 vccd1
+ vccd1 _22462_/A sky130_fd_sc_hd__mux4_1
XFILLER_33_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21412_ _21477_/A vssd1 vssd1 vccd1 vccd1 _21412_/X sky130_fd_sc_hd__clkbuf_1
X_24200_ _27572_/Q _24279_/A vssd1 vssd1 vccd1 vccd1 _24201_/A sky130_fd_sc_hd__and2_1
X_25180_ _25170_/A _25173_/B _25169_/Y vssd1 vssd1 vccd1 vccd1 _25181_/B sky130_fd_sc_hd__o21a_1
X_22392_ _22392_/A vssd1 vssd1 vccd1 vccd1 _22392_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24131_ _24175_/A vssd1 vssd1 vccd1 vccd1 _24140_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_175_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21343_ _21391_/A vssd1 vssd1 vccd1 vccd1 _21343_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1061 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24062_ _24062_/A vssd1 vssd1 vccd1 vccd1 _27308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21274_ _21290_/A vssd1 vssd1 vccd1 vccd1 _21274_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23013_ _23029_/A vssd1 vssd1 vccd1 vccd1 _23013_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20225_ _20225_/A vssd1 vssd1 vccd1 vccd1 _20225_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27821_ _25720_/X _27821_/D vssd1 vssd1 vccd1 vccd1 _27821_/Q sky130_fd_sc_hd__dfxtp_1
X_20156_ _20146_/X _20147_/X _20148_/X _20149_/X _20150_/X _20151_/X vssd1 vssd1 vccd1
+ vccd1 _20157_/A sky130_fd_sc_hd__mux4_1
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27752_ _27752_/CLK _27752_/D vssd1 vssd1 vccd1 vccd1 _27752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24964_ _24965_/A _24965_/B vssd1 vssd1 vccd1 vccd1 _24969_/B sky130_fd_sc_hd__nand2_1
X_20087_ _20087_/A vssd1 vssd1 vccd1 vccd1 _20087_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26703_ _21774_/X _26703_/D vssd1 vssd1 vccd1 vccd1 _26703_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23915_ _23913_/X _23914_/X _23938_/S vssd1 vssd1 vccd1 vccd1 _23915_/X sky130_fd_sc_hd__mux2_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27683_ _27791_/CLK _27683_/D vssd1 vssd1 vccd1 vccd1 _27974_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24895_ _27655_/Q _24885_/X _24894_/Y _24890_/X vssd1 vssd1 vccd1 vccd1 _27655_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26634_ _21528_/X _26634_/D vssd1 vssd1 vccd1 vccd1 _26634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23846_ _23844_/X _23845_/X _23846_/S vssd1 vssd1 vccd1 vccd1 _23846_/X sky130_fd_sc_hd__mux2_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26565_ _21292_/X _26565_/D vssd1 vssd1 vccd1 vccd1 _26565_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20989_ _20972_/X _20974_/X _20976_/X _20978_/X _20979_/X _20980_/X vssd1 vssd1 vccd1
+ vccd1 _20990_/A sky130_fd_sc_hd__mux4_1
X_23777_ _23777_/A vssd1 vssd1 vccd1 vccd1 _23777_/X sky130_fd_sc_hd__buf_2
XFILLER_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25516_ _27703_/Q _25509_/X _25510_/X vssd1 vssd1 vccd1 vccd1 _25516_/Y sky130_fd_sc_hd__a21oi_1
X_13530_ _13530_/A vssd1 vssd1 vccd1 vccd1 _13530_/X sky130_fd_sc_hd__buf_4
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22728_ _22728_/A vssd1 vssd1 vccd1 vccd1 _22728_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26496_ _21050_/X _26496_/D vssd1 vssd1 vccd1 vccd1 _26496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13461_ _26964_/Q _13435_/X _13457_/X _13460_/Y vssd1 vssd1 vccd1 vccd1 _26964_/D
+ sky130_fd_sc_hd__a31o_1
X_25447_ _24733_/A _25431_/X _25436_/Y _25444_/X _25446_/X vssd1 vssd1 vccd1 vccd1
+ _27755_/D sky130_fd_sc_hd__a221oi_1
X_22659_ _22649_/X _22650_/X _22651_/X _22652_/X _22653_/X _22654_/X vssd1 vssd1 vccd1
+ vccd1 _22660_/A sky130_fd_sc_hd__mux4_1
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15200_ _15200_/A vssd1 vssd1 vccd1 vccd1 _26358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16180_ _27576_/Q vssd1 vssd1 vccd1 vccd1 _16180_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13392_ _16235_/A vssd1 vssd1 vccd1 vccd1 _13392_/X sky130_fd_sc_hd__clkbuf_4
X_25378_ _27729_/Q input71/X _25380_/S vssd1 vssd1 vccd1 vccd1 _25379_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27117_ _27214_/CLK _27117_/D vssd1 vssd1 vccd1 vccd1 _27117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _15188_/S vssd1 vssd1 vccd1 vccd1 _15140_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24329_ _24329_/A vssd1 vssd1 vccd1 vccd1 _27448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27048_ _22970_/X _27048_/D vssd1 vssd1 vccd1 vccd1 _27048_/Q sky130_fd_sc_hd__dfxtp_1
X_15062_ _14731_/X _26419_/Q _15068_/S vssd1 vssd1 vccd1 vccd1 _15063_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14013_ _14032_/A vssd1 vssd1 vccd1 vccd1 _14029_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ _19886_/A vssd1 vssd1 vccd1 vccd1 _19870_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18821_ _19387_/A vssd1 vssd1 vccd1 vccd1 _18821_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18752_ _18752_/A vssd1 vssd1 vccd1 vccd1 _26036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15964_ _15967_/A vssd1 vssd1 vccd1 vccd1 _15964_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17703_ _25920_/Q _17702_/X _17706_/S vssd1 vssd1 vccd1 vccd1 _17704_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14915_ _14915_/A vssd1 vssd1 vccd1 vccd1 _26477_/D sky130_fd_sc_hd__clkbuf_1
X_18683_ _26006_/Q _17766_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _18684_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15895_ _15899_/A vssd1 vssd1 vccd1 vccd1 _15895_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17634_ _17469_/X _25889_/Q _17634_/S vssd1 vssd1 vccd1 vccd1 _17635_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14846_ _26507_/Q _13366_/X _14846_/S vssd1 vssd1 vccd1 vccd1 _14847_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _17472_/X _25858_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17566_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ _14775_/X _26533_/Q _14789_/S vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19304_ _19438_/A _19304_/B vssd1 vssd1 vccd1 vccd1 _19304_/X sky130_fd_sc_hd__or2_1
X_16516_ _25966_/Q _16311_/X _16515_/X vssd1 vssd1 vccd1 vccd1 _16805_/B sky130_fd_sc_hd__a21oi_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13728_ _13908_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13728_/Y sky130_fd_sc_hd__nor2_1
XFILLER_189_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17496_ _17495_/X _25833_/Q _17502_/S vssd1 vssd1 vccd1 vccd1 _17497_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19235_ _19226_/X _19230_/X _19234_/X _19186_/X _19139_/X vssd1 vssd1 vccd1 vccd1
+ _19246_/B sky130_fd_sc_hd__a221o_1
XFILLER_32_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16447_ _16722_/A _16447_/B _16447_/C _16447_/D vssd1 vssd1 vccd1 vccd1 _16447_/Y
+ sky130_fd_sc_hd__nor4_2
X_13659_ _13928_/A _13661_/B vssd1 vssd1 vccd1 vccd1 _13659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ _26151_/Q _26087_/Q _27015_/Q _26983_/Q _19165_/X _19070_/X vssd1 vssd1 vccd1
+ vccd1 _19167_/B sky130_fd_sc_hd__mux4_1
XFILLER_129_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16378_ _16378_/A vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18117_ _18392_/A vssd1 vssd1 vccd1 vccd1 _18117_/X sky130_fd_sc_hd__buf_2
X_15329_ _15329_/A vssd1 vssd1 vccd1 vccd1 _26300_/D sky130_fd_sc_hd__clkbuf_1
X_19097_ _19123_/A _19097_/B vssd1 vssd1 vccd1 vccd1 _19097_/X sky130_fd_sc_hd__or2_1
XFILLER_184_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18048_ _18305_/A vssd1 vssd1 vccd1 vccd1 _18048_/X sky130_fd_sc_hd__buf_2
XFILLER_99_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20010_ _20268_/A vssd1 vssd1 vccd1 vccd1 _20077_/A sky130_fd_sc_hd__buf_2
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19999_ _19999_/A vssd1 vssd1 vccd1 vccd1 _19999_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21961_ _21949_/X _21950_/X _21951_/X _21952_/X _21953_/X _21954_/X vssd1 vssd1 vccd1
+ vccd1 _21962_/A sky130_fd_sc_hd__mux4_1
XFILLER_95_993 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23700_ _23700_/A vssd1 vssd1 vccd1 vccd1 _27254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20912_ _20912_/A vssd1 vssd1 vccd1 vccd1 _20912_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21892_ _21892_/A vssd1 vssd1 vccd1 vccd1 _21892_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24680_ _27589_/Q _24673_/X _24679_/X _24677_/X vssd1 vssd1 vccd1 vccd1 _27589_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23631_ _25018_/A vssd1 vssd1 vccd1 vccd1 _25102_/S sky130_fd_sc_hd__buf_2
X_20843_ _20843_/A vssd1 vssd1 vccd1 vccd1 _20843_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26350_ _20541_/X _26350_/D vssd1 vssd1 vccd1 vccd1 _26350_/Q sky130_fd_sc_hd__dfxtp_1
X_23562_ _23562_/A vssd1 vssd1 vccd1 vccd1 _23577_/A sky130_fd_sc_hd__clkbuf_1
X_20774_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20852_/A sky130_fd_sc_hd__buf_2
XFILLER_161_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25301_ _25273_/A _25282_/A _25299_/Y _25295_/A _25300_/X vssd1 vssd1 vccd1 vccd1
+ _25329_/A sky130_fd_sc_hd__a41oi_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22513_ _22503_/X _22504_/X _22505_/X _22506_/X _22507_/X _22508_/X vssd1 vssd1 vccd1
+ vccd1 _22514_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23493_ _27190_/Q _23495_/B vssd1 vssd1 vccd1 vccd1 _23493_/X sky130_fd_sc_hd__or2_1
X_26281_ _20295_/X _26281_/D vssd1 vssd1 vccd1 vccd1 _26281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_28020_ _28020_/A _15983_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22444_ _22444_/A vssd1 vssd1 vccd1 vccd1 _22444_/X sky130_fd_sc_hd__clkbuf_1
X_25232_ _25229_/A _25228_/B _25228_/A vssd1 vssd1 vccd1 vccd1 _25266_/B sky130_fd_sc_hd__a21boi_2
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22375_ _22366_/X _22368_/X _22370_/X _22372_/X _22373_/X _22374_/X vssd1 vssd1 vccd1
+ vccd1 _22376_/A sky130_fd_sc_hd__mux4_1
X_25163_ _25149_/A _25146_/X _25149_/B _25155_/A _25147_/A vssd1 vssd1 vccd1 vccd1
+ _25164_/B sky130_fd_sc_hd__a311oi_2
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21326_ _21391_/A vssd1 vssd1 vccd1 vccd1 _21326_/X sky130_fd_sc_hd__clkbuf_1
X_24114_ _24114_/A vssd1 vssd1 vccd1 vccd1 _27331_/D sky130_fd_sc_hd__clkbuf_1
X_25094_ _25092_/X _25093_/X _27231_/Q vssd1 vssd1 vccd1 vccd1 _25094_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21257_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21257_/X sky130_fd_sc_hd__clkbuf_2
X_24045_ _24043_/X _24044_/X _24045_/S vssd1 vssd1 vccd1 vccd1 _24045_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20208_ _20200_/X _20201_/X _20202_/X _20203_/X _20204_/X _20205_/X vssd1 vssd1 vccd1
+ vccd1 _20209_/A sky130_fd_sc_hd__mux4_1
X_21188_ _21188_/A vssd1 vssd1 vccd1 vccd1 _21188_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27804_ _25668_/X _27804_/D vssd1 vssd1 vccd1 vccd1 _27804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20139_ _20139_/A vssd1 vssd1 vccd1 vccd1 _20139_/X sky130_fd_sc_hd__clkbuf_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25996_ _25996_/CLK _25996_/D vssd1 vssd1 vccd1 vccd1 _25996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27735_ _27735_/CLK _27735_/D vssd1 vssd1 vccd1 vccd1 _27735_/Q sky130_fd_sc_hd__dfxtp_1
X_12961_ _27816_/Q _12965_/B vssd1 vssd1 vccd1 vccd1 _12962_/A sky130_fd_sc_hd__and2_1
X_24947_ _24947_/A _24947_/B vssd1 vssd1 vccd1 vccd1 _24948_/B sky130_fd_sc_hd__nor2_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _26558_/Q _14698_/X _14693_/X _14699_/Y vssd1 vssd1 vccd1 vccd1 _26558_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27666_ _27666_/CLK _27666_/D vssd1 vssd1 vccd1 vccd1 _27666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15680_ _15680_/A vssd1 vssd1 vccd1 vccd1 _15689_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 _20607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24878_ _24889_/A _24878_/B vssd1 vssd1 vccd1 vccd1 _24878_/Y sky130_fd_sc_hd__nand2_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_311 _18152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 _19117_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26617_ _21470_/X _26617_/D vssd1 vssd1 vccd1 vccd1 _26617_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _15703_/A _14631_/B vssd1 vssd1 vccd1 vccd1 _14631_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_333 _13111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23829_ _23827_/X _23828_/X _23844_/S vssd1 vssd1 vccd1 vccd1 _23829_/X sky130_fd_sc_hd__mux2_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_344 _13389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27597_ _27597_/CLK _27597_/D vssd1 vssd1 vccd1 vccd1 _27597_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 _14718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_366 _26814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _25940_/Q _26006_/Q _17370_/S vssd1 vssd1 vccd1 vccd1 _17351_/B sky130_fd_sc_hd__mux2_1
XANTENNA_377 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _26609_/Q _14549_/X _14553_/X _14561_/Y vssd1 vssd1 vccd1 vccd1 _26609_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26548_ _21226_/X _26548_/D vssd1 vssd1 vccd1 vccd1 _26548_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16301_ _16798_/A _16301_/B _16301_/C _16301_/D vssd1 vssd1 vccd1 vccd1 _16576_/B
+ sky130_fd_sc_hd__or4_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13902_/A _13517_/B vssd1 vssd1 vccd1 vccd1 _13513_/Y sky130_fd_sc_hd__nor2_1
X_17281_ input37/X vssd1 vssd1 vccd1 vccd1 _17281_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14493_/A vssd1 vssd1 vccd1 vccd1 _15754_/A sky130_fd_sc_hd__clkbuf_2
X_26479_ _20990_/X _26479_/D vssd1 vssd1 vccd1 vccd1 _26479_/Q sky130_fd_sc_hd__dfxtp_1
X_19020_ _27800_/Q _26561_/Q _26433_/Q _26113_/Q _18974_/X _19019_/X vssd1 vssd1 vccd1
+ vccd1 _19020_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16232_ _15992_/A _16228_/X _16229_/X _16230_/X _16231_/X vssd1 vssd1 vccd1 vccd1
+ _16408_/A sky130_fd_sc_hd__o41a_1
X_13444_ _27363_/Q _13019_/A _13027_/A _27331_/Q _13070_/X vssd1 vssd1 vccd1 vccd1
+ _16134_/A sky130_fd_sc_hd__a221oi_4
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16163_ _26053_/Q _16274_/B _16298_/C vssd1 vssd1 vccd1 vccd1 _16445_/B sky130_fd_sc_hd__and3_1
X_13375_ _13375_/A vssd1 vssd1 vccd1 vccd1 _26985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ _14807_/X _26395_/Q _15116_/S vssd1 vssd1 vccd1 vccd1 _15115_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16094_ _16094_/A vssd1 vssd1 vccd1 vccd1 _16094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19922_ _25657_/A vssd1 vssd1 vccd1 vccd1 _20270_/A sky130_fd_sc_hd__clkbuf_1
X_15045_ _15334_/B _15045_/B _15334_/C vssd1 vssd1 vccd1 vccd1 _15262_/B sky130_fd_sc_hd__nand3b_4
XFILLER_141_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19853_ _19901_/A vssd1 vssd1 vccd1 vccd1 _19853_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18804_ _19296_/S vssd1 vssd1 vccd1 vccd1 _19299_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_394 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19784_ _19800_/A vssd1 vssd1 vccd1 vccd1 _19784_/X sky130_fd_sc_hd__clkbuf_2
X_16996_ _16992_/X _16996_/B vssd1 vssd1 vccd1 vccd1 _16996_/X sky130_fd_sc_hd__and2b_1
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18735_ _26029_/Q _17737_/X _18735_/S vssd1 vssd1 vccd1 vccd1 _18736_/A sky130_fd_sc_hd__mux2_1
X_15947_ _15949_/A vssd1 vssd1 vccd1 vccd1 _15947_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18666_ _25998_/Q _17740_/X _18674_/S vssd1 vssd1 vccd1 vccd1 _18667_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _15881_/A vssd1 vssd1 vccd1 vccd1 _15878_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14829_ _26515_/Q _13341_/X _14835_/S vssd1 vssd1 vccd1 vccd1 _14830_/A sky130_fd_sc_hd__mux2_1
X_17617_ _17444_/X _25881_/Q _17623_/S vssd1 vssd1 vccd1 vccd1 _17618_/A sky130_fd_sc_hd__mux2_1
X_18597_ _27540_/Q _27519_/Q vssd1 vssd1 vccd1 vccd1 _18598_/B sky130_fd_sc_hd__or2_1
XFILLER_184_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17548_ _17548_/A vssd1 vssd1 vccd1 vccd1 _25850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17479_ _27425_/Q vssd1 vssd1 vccd1 vccd1 _17479_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19218_ _26281_/Q _26249_/Q _26217_/Q _26185_/Q _18778_/X _18782_/X vssd1 vssd1 vccd1
+ vccd1 _19218_/X sky130_fd_sc_hd__mux4_2
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20490_ _20480_/X _20481_/X _20482_/X _20483_/X _20484_/X _20485_/X vssd1 vssd1 vccd1
+ vccd1 _20491_/A sky130_fd_sc_hd__mux4_1
XFILLER_9_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19149_ _26534_/Q _26502_/Q _26470_/Q _27046_/Q _19102_/X _19148_/X vssd1 vssd1 vccd1
+ vccd1 _19149_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22160_ _22176_/A vssd1 vssd1 vccd1 vccd1 _22160_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21111_ _21127_/A vssd1 vssd1 vccd1 vccd1 _21111_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22091_ _22083_/X _22084_/X _22085_/X _22086_/X _22088_/X _22090_/X vssd1 vssd1 vccd1
+ vccd1 _22092_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21042_ _21042_/A vssd1 vssd1 vccd1 vccd1 _21042_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25850_ _25985_/CLK _25850_/D vssd1 vssd1 vccd1 vccd1 _25850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24801_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24801_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25781_ _25792_/A vssd1 vssd1 vccd1 vccd1 _25790_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22993_ _25635_/A vssd1 vssd1 vccd1 vccd1 _22993_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27520_ _27520_/CLK _27520_/D vssd1 vssd1 vccd1 vccd1 _27520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24732_ _24554_/A _24727_/X _24731_/X _24729_/X vssd1 vssd1 vccd1 vccd1 _27609_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21944_ _21944_/A vssd1 vssd1 vccd1 vccd1 _21944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27985__451 vssd1 vssd1 vccd1 vccd1 _27985__451/HI _27985_/A sky130_fd_sc_hd__conb_1
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27451_ _27454_/CLK _27451_/D vssd1 vssd1 vccd1 vccd1 _27451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24663_ _24663_/A vssd1 vssd1 vccd1 vccd1 _24663_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21875_ _21863_/X _21864_/X _21865_/X _21866_/X _21867_/X _21868_/X vssd1 vssd1 vccd1
+ vccd1 _21876_/A sky130_fd_sc_hd__mux4_1
XFILLER_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26402_ _20717_/X _26402_/D vssd1 vssd1 vccd1 vccd1 _26402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23614_ _23614_/A vssd1 vssd1 vccd1 vccd1 _27223_/D sky130_fd_sc_hd__clkbuf_1
X_20826_ _20816_/X _20817_/X _20818_/X _20819_/X _20820_/X _20821_/X vssd1 vssd1 vccd1
+ vccd1 _20827_/A sky130_fd_sc_hd__mux4_1
X_27382_ _27407_/CLK _27382_/D vssd1 vssd1 vccd1 vccd1 _27382_/Q sky130_fd_sc_hd__dfxtp_1
X_24594_ _27657_/Q _24598_/B vssd1 vssd1 vccd1 vccd1 _24595_/A sky130_fd_sc_hd__and2_1
XFILLER_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26333_ _20477_/X _26333_/D vssd1 vssd1 vccd1 vccd1 _26333_/Q sky130_fd_sc_hd__dfxtp_1
X_23545_ _23562_/A vssd1 vssd1 vccd1 vccd1 _23560_/A sky130_fd_sc_hd__clkbuf_1
X_20757_ _20773_/A vssd1 vssd1 vccd1 vccd1 _20757_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26264_ _20231_/X _26264_/D vssd1 vssd1 vccd1 vccd1 _26264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_898 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20688_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20758_/A sky130_fd_sc_hd__clkbuf_2
X_23476_ _27183_/Q _23483_/B vssd1 vssd1 vccd1 vccd1 _23476_/X sky130_fd_sc_hd__or2_1
XFILLER_10_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_28003_ _28003_/A _15877_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_25215_ _27702_/Q _25184_/X _25213_/Y _25214_/X vssd1 vssd1 vccd1 vccd1 _27702_/D
+ sky130_fd_sc_hd__o211a_1
X_22427_ _22417_/X _22418_/X _22419_/X _22420_/X _22421_/X _22422_/X vssd1 vssd1 vccd1
+ vccd1 _22428_/A sky130_fd_sc_hd__mux4_1
XFILLER_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26195_ _19999_/X _26195_/D vssd1 vssd1 vccd1 vccd1 _26195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25146_ _27524_/Q _27492_/Q vssd1 vssd1 vccd1 vccd1 _25146_/X sky130_fd_sc_hd__or2_1
XFILLER_108_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13160_ _27348_/Q _13021_/A _13102_/X _27316_/Q _13159_/X vssd1 vssd1 vccd1 vccd1
+ _14769_/A sky130_fd_sc_hd__a221o_4
XFILLER_200_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22358_ _22358_/A vssd1 vssd1 vccd1 vccd1 _22358_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21309_ _21653_/A vssd1 vssd1 vccd1 vccd1 _21378_/A sky130_fd_sc_hd__clkbuf_2
X_13091_ _13530_/A vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__clkbuf_2
X_22289_ _22280_/X _22282_/X _22284_/X _22286_/X _22287_/X _22288_/X vssd1 vssd1 vccd1
+ vccd1 _22290_/A sky130_fd_sc_hd__mux4_1
X_25077_ _25077_/A vssd1 vssd1 vccd1 vccd1 _27683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27953__439 vssd1 vssd1 vccd1 vccd1 _27953__439/HI _27953_/A sky130_fd_sc_hd__conb_1
XFILLER_85_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24028_ _23990_/X _24026_/X _24027_/X _24005_/X vssd1 vssd1 vccd1 vccd1 _27299_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16850_ _16841_/X _16844_/X _16846_/Y _16849_/X vssd1 vssd1 vccd1 vccd1 _24215_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15801_ _13099_/X _26098_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15802_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16781_ _16779_/Y _16780_/X _16770_/Y vssd1 vssd1 vccd1 vccd1 _16781_/X sky130_fd_sc_hd__a21o_1
X_13993_ _26797_/Q _13987_/X _13983_/X _13992_/Y vssd1 vssd1 vccd1 vccd1 _26797_/D
+ sky130_fd_sc_hd__a31o_1
X_25979_ _26018_/CLK _25979_/D vssd1 vssd1 vccd1 vccd1 _25979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18520_ _26550_/Q _26518_/Q _26486_/Q _27062_/Q _17999_/X _17901_/X vssd1 vssd1 vccd1
+ vccd1 _18520_/X sky130_fd_sc_hd__mux4_1
X_15732_ _15732_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15732_/Y sky130_fd_sc_hd__nor2_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27718_ _27719_/CLK _27718_/D vssd1 vssd1 vccd1 vccd1 _27718_/Q sky130_fd_sc_hd__dfxtp_1
X_12944_ _27823_/Q _12952_/B vssd1 vssd1 vccd1 vccd1 _12945_/A sky130_fd_sc_hd__and2_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _18451_/A _17910_/X vssd1 vssd1 vccd1 vccd1 _18451_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27649_ _27649_/CLK _27649_/D vssd1 vssd1 vccd1 vccd1 _27649_/Q sky130_fd_sc_hd__dfxtp_1
X_15663_ _13156_/X _26152_/Q _15667_/S vssd1 vssd1 vccd1 vccd1 _15664_/A sky130_fd_sc_hd__mux2_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _23946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _25106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _13198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17402_ _25639_/A vssd1 vssd1 vccd1 vccd1 _19625_/A sky130_fd_sc_hd__buf_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _25106_/A vssd1 vssd1 vccd1 vccd1 _14671_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _26704_/Q _26672_/Q _26640_/Q _26608_/Q _18360_/X _18249_/X vssd1 vssd1 vccd1
+ vccd1 _18383_/A sky130_fd_sc_hd__mux4_2
XANTENNA_163 _13385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15594_ _15594_/A vssd1 vssd1 vccd1 vccd1 _26183_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _14471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 _16442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17333_ _27092_/Q _27124_/Q _17355_/S vssd1 vssd1 vccd1 vccd1 _17333_/X sky130_fd_sc_hd__mux2_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14558_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17264_ _17325_/A vssd1 vssd1 vccd1 vccd1 _17264_/X sky130_fd_sc_hd__buf_2
XFILLER_144_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ _15741_/A _14483_/B vssd1 vssd1 vccd1 vccd1 _14476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19003_ _26144_/Q _26080_/Q _27008_/Q _26976_/Q _18882_/X _18950_/X vssd1 vssd1 vccd1
+ vccd1 _19004_/B sky130_fd_sc_hd__mux4_1
X_16215_ _26046_/Q _16215_/B _16221_/C vssd1 vssd1 vccd1 vccd1 _16215_/X sky130_fd_sc_hd__and3_1
X_13427_ _13762_/B _15335_/A vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__or2_1
X_17195_ _25826_/Q _26025_/Q _17219_/S vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16146_ _16110_/A _24302_/A _16623_/A vssd1 vssd1 vccd1 vccd1 _16797_/A sky130_fd_sc_hd__o21ai_1
X_13358_ _26990_/Q _13357_/X _13367_/S vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16077_ _16077_/A vssd1 vssd1 vccd1 vccd1 _16077_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289_ _27015_/Q _13161_/X _13291_/S vssd1 vssd1 vccd1 vccd1 _13290_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15028_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15028_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19905_ _19977_/A vssd1 vssd1 vccd1 vccd1 _19905_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19836_ _19836_/A vssd1 vssd1 vccd1 vccd1 _19901_/A sky130_fd_sc_hd__buf_2
XFILLER_190_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19767_ _19815_/A vssd1 vssd1 vccd1 vccd1 _19767_/X sky130_fd_sc_hd__clkbuf_1
X_16979_ _16979_/A _16979_/B _27590_/Q vssd1 vssd1 vccd1 vccd1 _16980_/C sky130_fd_sc_hd__and3_1
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18718_ _26021_/Q _17712_/X _18724_/S vssd1 vssd1 vccd1 vccd1 _18719_/A sky130_fd_sc_hd__mux2_1
X_19698_ _19714_/A vssd1 vssd1 vccd1 vccd1 _19698_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_462 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18649_ _18649_/A vssd1 vssd1 vccd1 vccd1 _25990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21660_ _21660_/A vssd1 vssd1 vccd1 vccd1 _21660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20611_ _20611_/A vssd1 vssd1 vccd1 vccd1 _20611_/X sky130_fd_sc_hd__clkbuf_1
X_21591_ _21580_/X _21582_/X _21584_/X _21586_/X _21587_/X _21588_/X vssd1 vssd1 vccd1
+ vccd1 _21592_/A sky130_fd_sc_hd__mux4_1
X_23330_ input53/X input54/X input55/X input56/X vssd1 vssd1 vccd1 vccd1 _23331_/D
+ sky130_fd_sc_hd__or4_1
X_20542_ _20531_/X _20533_/X _20535_/X _20537_/X _20538_/X _20539_/X vssd1 vssd1 vccd1
+ vccd1 _20543_/A sky130_fd_sc_hd__mux4_1
XFILLER_193_824 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20473_ _20473_/A vssd1 vssd1 vccd1 vccd1 _20473_/X sky130_fd_sc_hd__clkbuf_1
X_23261_ input60/X vssd1 vssd1 vccd1 vccd1 _23261_/Y sky130_fd_sc_hd__inv_2
X_25000_ _25000_/A vssd1 vssd1 vccd1 vccd1 _27674_/D sky130_fd_sc_hd__clkbuf_1
X_22212_ _22212_/A vssd1 vssd1 vccd1 vccd1 _22212_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23192_ _23192_/A vssd1 vssd1 vccd1 vccd1 _27133_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22143_ _22175_/A vssd1 vssd1 vccd1 vccd1 _22143_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22074_ _22074_/A vssd1 vssd1 vccd1 vccd1 _22074_/X sky130_fd_sc_hd__clkbuf_1
X_26951_ _22642_/X _26951_/D vssd1 vssd1 vccd1 vccd1 _26951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25902_ _27157_/CLK _25902_/D vssd1 vssd1 vccd1 vccd1 _25902_/Q sky130_fd_sc_hd__dfxtp_1
X_21025_ _21041_/A vssd1 vssd1 vccd1 vccd1 _21025_/X sky130_fd_sc_hd__clkbuf_1
X_26882_ _22396_/X _26882_/D vssd1 vssd1 vccd1 vccd1 _26882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25833_ _27151_/CLK _25833_/D vssd1 vssd1 vccd1 vccd1 _25833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25764_ _17463_/X _27838_/Q _25768_/S vssd1 vssd1 vccd1 vccd1 _25765_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22976_ _25636_/A vssd1 vssd1 vccd1 vccd1 _22976_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27503_ _27627_/CLK _27503_/D vssd1 vssd1 vccd1 vccd1 _27503_/Q sky130_fd_sc_hd__dfxtp_1
X_24715_ _25434_/A vssd1 vssd1 vccd1 vccd1 _24725_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_71_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21927_ _21911_/X _21912_/X _21913_/X _21914_/X _21916_/X _21918_/X vssd1 vssd1 vccd1
+ vccd1 _21928_/A sky130_fd_sc_hd__mux4_1
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25695_ _25689_/X _25690_/X _25691_/X _25692_/X _25693_/X _25694_/X vssd1 vssd1 vccd1
+ vccd1 _25696_/A sky130_fd_sc_hd__mux4_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27434_ _27435_/CLK _27434_/D vssd1 vssd1 vccd1 vccd1 _27434_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24646_ _27162_/Q _24658_/B vssd1 vssd1 vccd1 vccd1 _24646_/X sky130_fd_sc_hd__or2_1
X_21858_ _21858_/A vssd1 vssd1 vccd1 vccd1 _21858_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20809_/A vssd1 vssd1 vccd1 vccd1 _20809_/X sky130_fd_sc_hd__clkbuf_1
X_27365_ _27365_/CLK _27365_/D vssd1 vssd1 vccd1 vccd1 _27365_/Q sky130_fd_sc_hd__dfxtp_1
X_24577_ _24577_/A vssd1 vssd1 vccd1 vccd1 _27549_/D sky130_fd_sc_hd__clkbuf_1
X_21789_ _21777_/X _21778_/X _21779_/X _21780_/X _21781_/X _21782_/X vssd1 vssd1 vccd1
+ vccd1 _21790_/A sky130_fd_sc_hd__mux4_1
XFILLER_196_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14330_ _14344_/A vssd1 vssd1 vccd1 vccd1 _14335_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_26316_ _20417_/X _26316_/D vssd1 vssd1 vccd1 vccd1 _26316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23528_ _23562_/A vssd1 vssd1 vccd1 vccd1 _23543_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_27296_ _27296_/CLK _27296_/D vssd1 vssd1 vccd1 vccd1 _27296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14261_ _14348_/A _14263_/B vssd1 vssd1 vccd1 vccd1 _14261_/Y sky130_fd_sc_hd__nor2_1
X_26247_ _20175_/X _26247_/D vssd1 vssd1 vccd1 vccd1 _26247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23459_ _27177_/Q _23470_/B vssd1 vssd1 vccd1 vccd1 _23459_/X sky130_fd_sc_hd__or2_1
XFILLER_125_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16000_ _27480_/Q _27371_/Q vssd1 vssd1 vccd1 vccd1 _16001_/D sky130_fd_sc_hd__xnor2_1
XFILLER_143_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ _13212_/A vssd1 vssd1 vccd1 vccd1 _27039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14192_ _14369_/A _14200_/B vssd1 vssd1 vccd1 vccd1 _14192_/Y sky130_fd_sc_hd__nor2_1
X_26178_ _19937_/X _26178_/D vssd1 vssd1 vccd1 vccd1 _26178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25129_ _25129_/A _25129_/B vssd1 vssd1 vccd1 vccd1 _25130_/B sky130_fd_sc_hd__nand2_1
X_13143_ _27351_/Q _13090_/X _13091_/X _27319_/Q _13142_/X vssd1 vssd1 vccd1 vccd1
+ _14759_/A sky130_fd_sc_hd__a221o_4
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _18425_/A vssd1 vssd1 vccd1 vccd1 _17951_/X sky130_fd_sc_hd__clkbuf_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _13074_/A vssd1 vssd1 vccd1 vccd1 _27062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16902_ _16902_/A _16902_/B vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__nor2_1
X_17882_ _17882_/A vssd1 vssd1 vccd1 vccd1 _25945_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater309 _27467_/CLK vssd1 vssd1 vccd1 vccd1 _27468_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_120_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19621_ _19637_/A vssd1 vssd1 vccd1 vccd1 _19621_/X sky130_fd_sc_hd__clkbuf_1
X_16833_ _16833_/A _16916_/A vssd1 vssd1 vccd1 vccd1 _16833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19552_ _27824_/Q _26585_/Q _26457_/Q _26137_/Q _18922_/X _18923_/X vssd1 vssd1 vccd1
+ vccd1 _19552_/X sky130_fd_sc_hd__mux4_1
X_16764_ _16764_/A _16764_/B vssd1 vssd1 vccd1 vccd1 _16765_/C sky130_fd_sc_hd__xor2_1
X_13976_ _14448_/A vssd1 vssd1 vccd1 vccd1 _14354_/A sky130_fd_sc_hd__buf_2
X_15715_ _26132_/Q _15705_/X _15713_/X _15714_/Y vssd1 vssd1 vccd1 vccd1 _26132_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18503_ _26293_/Q _26261_/Q _26229_/Q _26197_/Q _18458_/X _18481_/X vssd1 vssd1 vccd1
+ vccd1 _18503_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12927_ input48/X input49/X input50/X input51/X vssd1 vssd1 vccd1 vccd1 _12928_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_20_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19483_ _26165_/Q _26101_/Q _27029_/Q _26997_/Q _19460_/X _19482_/X vssd1 vssd1 vccd1
+ vccd1 _19484_/B sky130_fd_sc_hd__mux4_1
X_16695_ _16619_/X _16609_/B _16692_/X _16694_/X vssd1 vssd1 vccd1 vccd1 _24237_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_111_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18434_ _18311_/X _18429_/X _18433_/X _18412_/X vssd1 vssd1 vccd1 vccd1 _18445_/B
+ sky130_fd_sc_hd__a211o_1
X_15646_ _15646_/A vssd1 vssd1 vccd1 vccd1 _26160_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ _26543_/Q _26511_/Q _26479_/Q _27055_/Q _17899_/X _17901_/X vssd1 vssd1 vccd1
+ vccd1 _18365_/X sky130_fd_sc_hd__mux4_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15577_ _15577_/A vssd1 vssd1 vccd1 vccd1 _26191_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17277_/X _17316_/B vssd1 vssd1 vccd1 vccd1 _17316_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14528_ _15779_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14528_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18296_ _27597_/Q vssd1 vssd1 vccd1 vccd1 _18352_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_187_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _27085_/Q _27117_/Q _17295_/S vssd1 vssd1 vccd1 vccd1 _17247_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14459_ _14548_/A vssd1 vssd1 vccd1 vccd1 _14530_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17178_ _27840_/Q _27144_/Q _25889_/Q _25857_/Q _17142_/X _17130_/X vssd1 vssd1 vccd1
+ vccd1 _17178_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16129_ _16036_/X _24308_/A _16648_/A vssd1 vssd1 vccd1 vccd1 _16792_/A sky130_fd_sc_hd__o21a_1
XFILLER_6_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ _19887_/A vssd1 vssd1 vccd1 vccd1 _19819_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22830_ _22830_/A vssd1 vssd1 vccd1 vccd1 _22830_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22761_ _22751_/X _22752_/X _22753_/X _22754_/X _22755_/X _22756_/X vssd1 vssd1 vccd1
+ vccd1 _22762_/A sky130_fd_sc_hd__mux4_1
XFILLER_198_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24500_ _24400_/A _24633_/C _24498_/X _24499_/X vssd1 vssd1 vccd1 vccd1 _27520_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21712_ _21712_/A vssd1 vssd1 vccd1 vccd1 _21712_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25480_ _25569_/A vssd1 vssd1 vccd1 vccd1 _25480_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22692_ _22692_/A vssd1 vssd1 vccd1 vccd1 _22692_/X sky130_fd_sc_hd__clkbuf_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24431_ _27615_/Q _24433_/B vssd1 vssd1 vccd1 vccd1 _24432_/A sky130_fd_sc_hd__and2_1
X_21643_ _21631_/X _21632_/X _21633_/X _21634_/X _21635_/X _21636_/X vssd1 vssd1 vccd1
+ vccd1 _21644_/A sky130_fd_sc_hd__mux4_1
XFILLER_178_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27150_ _27154_/CLK _27150_/D vssd1 vssd1 vccd1 vccd1 _27150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24362_ _24362_/A vssd1 vssd1 vccd1 vccd1 _27463_/D sky130_fd_sc_hd__clkbuf_1
X_21574_ _21574_/A vssd1 vssd1 vccd1 vccd1 _21574_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_30 _27837_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _17810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_52 _18102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26101_ _19671_/X _26101_/D vssd1 vssd1 vccd1 vccd1 _26101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23313_ _27723_/Q _23281_/Y _23312_/Y input54/X vssd1 vssd1 vccd1 vccd1 _23313_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_63 _18307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27081_ _27081_/CLK _27081_/D vssd1 vssd1 vccd1 vccd1 _27081_/Q sky130_fd_sc_hd__dfxtp_1
X_20525_ _20525_/A vssd1 vssd1 vccd1 vccd1 _20525_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24293_ _24293_/A _24302_/B vssd1 vssd1 vccd1 vccd1 _27424_/D sky130_fd_sc_hd__nor2_1
XANTENNA_74 _18488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_85 _18930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 _19210_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26032_ _27151_/CLK _26032_/D vssd1 vssd1 vccd1 vccd1 _26032_/Q sky130_fd_sc_hd__dfxtp_1
X_23244_ _17511_/X _27157_/Q _23248_/S vssd1 vssd1 vccd1 vccd1 _23245_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20456_ _20445_/X _20447_/X _20449_/X _20451_/X _20452_/X _20453_/X vssd1 vssd1 vccd1
+ vccd1 _20457_/A sky130_fd_sc_hd__mux4_1
XFILLER_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23175_ _23175_/A vssd1 vssd1 vccd1 vccd1 _27126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20387_ _20387_/A vssd1 vssd1 vccd1 vccd1 _20387_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22126_ _22174_/A vssd1 vssd1 vccd1 vccd1 _22126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_701 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27983_ _27983_/A _15899_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
XFILLER_161_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26934_ _22576_/X _26934_/D vssd1 vssd1 vccd1 vccd1 _26934_/Q sky130_fd_sc_hd__dfxtp_1
X_22057_ _22051_/X _22052_/X _22053_/X _22054_/X _22055_/X _22056_/X vssd1 vssd1 vccd1
+ vccd1 _22058_/A sky130_fd_sc_hd__mux4_1
XFILLER_47_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21008_ _21040_/A vssd1 vssd1 vccd1 vccd1 _21008_/X sky130_fd_sc_hd__clkbuf_1
X_26865_ _22338_/X _26865_/D vssd1 vssd1 vccd1 vccd1 _26865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _13923_/A _13838_/B vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__nor2_1
X_25816_ _27414_/CLK _25816_/D vssd1 vssd1 vccd1 vccd1 _25816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26796_ _22094_/X _26796_/D vssd1 vssd1 vccd1 vccd1 _26796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13761_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13761_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25747_ _25747_/A vssd1 vssd1 vccd1 vccd1 _27830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22959_ _22959_/A vssd1 vssd1 vccd1 vccd1 _23029_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15500_ _15500_/A vssd1 vssd1 vccd1 vccd1 _26225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _16475_/Y _16890_/A _16433_/B _16719_/B _16479_/Y vssd1 vssd1 vccd1 vccd1
+ _16481_/A sky130_fd_sc_hd__o221a_1
X_13692_ _13745_/A vssd1 vssd1 vccd1 vccd1 _13692_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25678_ _25710_/A vssd1 vssd1 vccd1 vccd1 _25678_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27417_ _27417_/CLK _27417_/D vssd1 vssd1 vccd1 vccd1 _27417_/Q sky130_fd_sc_hd__dfxtp_1
X_15431_ _15477_/S vssd1 vssd1 vccd1 vccd1 _15440_/S sky130_fd_sc_hd__clkbuf_2
X_24629_ _24638_/A _24629_/B vssd1 vssd1 vccd1 vccd1 _24630_/A sky130_fd_sc_hd__and2_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18150_ _18150_/A vssd1 vssd1 vccd1 vccd1 _18150_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15362_ _14747_/X _26286_/Q _15368_/S vssd1 vssd1 vccd1 vccd1 _15363_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27348_ _27348_/CLK _27348_/D vssd1 vssd1 vccd1 vccd1 _27348_/Q sky130_fd_sc_hd__dfxtp_2
X_17101_ _27073_/Q _27105_/Q _17112_/S vssd1 vssd1 vccd1 vccd1 _17101_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14313_ _26688_/Q _14310_/X _14311_/X _14312_/Y vssd1 vssd1 vccd1 vccd1 _26688_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18081_ _18156_/A vssd1 vssd1 vccd1 vccd1 _18514_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15293_ _26316_/Q _13363_/X _15295_/S vssd1 vssd1 vccd1 vccd1 _15294_/A sky130_fd_sc_hd__mux2_1
X_27279_ _27308_/CLK _27279_/D vssd1 vssd1 vccd1 vccd1 _27279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27959__445 vssd1 vssd1 vccd1 vccd1 _27959__445/HI _27959_/A sky130_fd_sc_hd__conb_1
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17032_ _25813_/Q _26012_/Q _17061_/A vssd1 vssd1 vccd1 vccd1 _17032_/X sky130_fd_sc_hd__mux2_1
X_14244_ _14331_/A _14248_/B vssd1 vssd1 vccd1 vccd1 _14244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14175_ _26738_/Q _14173_/X _14167_/X _14174_/Y vssd1 vssd1 vccd1 vccd1 _26738_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _27354_/Q _13063_/A _13082_/X _27322_/Q _13125_/X vssd1 vssd1 vccd1 vccd1
+ _13127_/A sky130_fd_sc_hd__a221o_1
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18983_ _26399_/Q _26367_/Q _26335_/Q _26303_/Q _18887_/X _18982_/X vssd1 vssd1 vccd1
+ vccd1 _18983_/X sky130_fd_sc_hd__mux4_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _26141_/Q _26077_/Q _27005_/Q _26973_/Q _17870_/X _17824_/X vssd1 vssd1 vccd1
+ vccd1 _17936_/A sky130_fd_sc_hd__mux4_1
X_13057_ _27365_/Q _13022_/X _13030_/X _27333_/Q _13056_/X vssd1 vssd1 vccd1 vccd1
+ _14715_/A sky130_fd_sc_hd__a221o_1
XFILLER_87_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater106 _25900_/CLK vssd1 vssd1 vccd1 vccd1 _27851_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater117 _27684_/CLK vssd1 vssd1 vccd1 vccd1 _27214_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater128 _26038_/CLK vssd1 vssd1 vccd1 vccd1 _25941_/CLK sky130_fd_sc_hd__clkbuf_1
X_17865_ _18177_/A vssd1 vssd1 vccd1 vccd1 _17865_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater139 _26026_/CLK vssd1 vssd1 vccd1 vccd1 _27145_/CLK sky130_fd_sc_hd__clkbuf_1
X_19604_ _19604_/A vssd1 vssd1 vccd1 vccd1 _19604_/X sky130_fd_sc_hd__clkbuf_1
X_16816_ _16816_/A _16816_/B vssd1 vssd1 vccd1 vccd1 _16816_/Y sky130_fd_sc_hd__nand2_1
X_17796_ _17786_/X _17792_/X _17886_/S vssd1 vssd1 vccd1 vccd1 _17796_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19535_ _26712_/Q _26680_/Q _26648_/Q _26616_/Q _18816_/X _18818_/X vssd1 vssd1 vccd1
+ vccd1 _19535_/X sky130_fd_sc_hd__mux4_1
X_13959_ _14340_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _13959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16747_ _16747_/A _16747_/B vssd1 vssd1 vccd1 vccd1 _16765_/A sky130_fd_sc_hd__xor2_1
XFILLER_185_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19466_ _26420_/Q _26388_/Q _26356_/Q _26324_/Q _19465_/X _19399_/X vssd1 vssd1 vccd1
+ vccd1 _19466_/X sky130_fd_sc_hd__mux4_1
X_16678_ _16393_/Y _16738_/B _16715_/C vssd1 vssd1 vccd1 vccd1 _16678_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18417_ _18279_/X _18416_/X _18326_/X vssd1 vssd1 vccd1 vccd1 _18417_/X sky130_fd_sc_hd__o21a_1
X_15629_ _15629_/A vssd1 vssd1 vccd1 vccd1 _26168_/D sky130_fd_sc_hd__clkbuf_1
X_19397_ _26289_/Q _26257_/Q _26225_/Q _26193_/Q _19283_/X _19352_/X vssd1 vssd1 vccd1
+ vccd1 _19397_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18348_ _26542_/Q _26510_/Q _26478_/Q _27054_/Q _18011_/A _18141_/A vssd1 vssd1 vccd1
+ vccd1 _18348_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18279_ _18437_/A vssd1 vssd1 vccd1 vccd1 _18279_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20310_ _20302_/X _20303_/X _20304_/X _20305_/X _20306_/X _20307_/X vssd1 vssd1 vccd1
+ vccd1 _20311_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput50 la1_oenb[18] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_6
X_21290_ _21290_/A vssd1 vssd1 vccd1 vccd1 _21290_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 la1_oenb[28] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_4
Xinput72 la1_oenb[9] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_4
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20241_ _20241_/A vssd1 vssd1 vccd1 vccd1 _20241_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20172_ _20162_/X _20163_/X _20164_/X _20165_/X _20167_/X _20169_/X vssd1 vssd1 vccd1
+ vccd1 _20173_/A sky130_fd_sc_hd__mux4_1
XFILLER_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24980_ _27963_/A _24979_/X _24980_/S vssd1 vssd1 vccd1 vccd1 _24981_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23931_ _23928_/X _23930_/X _23938_/S vssd1 vssd1 vccd1 vccd1 _23931_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26650_ _21590_/X _26650_/D vssd1 vssd1 vccd1 vccd1 _26650_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23862_ _23862_/A vssd1 vssd1 vccd1 vccd1 _23862_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28010__476 vssd1 vssd1 vccd1 vccd1 _28010__476/HI _28010_/A sky130_fd_sc_hd__conb_1
XFILLER_26_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25601_ _25601_/A _25601_/B vssd1 vssd1 vccd1 vccd1 _25601_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22813_ _22802_/X _22804_/X _22806_/X _22808_/X _22809_/X _22810_/X vssd1 vssd1 vccd1
+ vccd1 _22814_/A sky130_fd_sc_hd__mux4_1
X_26581_ _21350_/X _26581_/D vssd1 vssd1 vccd1 vccd1 _26581_/Q sky130_fd_sc_hd__dfxtp_1
X_23793_ _27830_/Q _27134_/Q _25879_/Q _25847_/Q _23777_/X _23744_/X vssd1 vssd1 vccd1
+ vccd1 _23793_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25532_ _25530_/X _25237_/B _25531_/X _25513_/X vssd1 vssd1 vccd1 vccd1 _25532_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22744_ _22744_/A vssd1 vssd1 vccd1 vccd1 _22744_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25463_ _25524_/A vssd1 vssd1 vccd1 vccd1 _25463_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22675_ _22665_/X _22666_/X _22667_/X _22668_/X _22669_/X _22670_/X vssd1 vssd1 vccd1
+ vccd1 _22676_/A sky130_fd_sc_hd__mux4_1
XFILLER_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27202_ _27208_/CLK _27202_/D vssd1 vssd1 vccd1 vccd1 _27202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24414_ _27587_/Q _24422_/B vssd1 vssd1 vccd1 vccd1 _24415_/A sky130_fd_sc_hd__and2_1
X_21626_ _21626_/A vssd1 vssd1 vccd1 vccd1 _21626_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25394_ _27736_/Q input47/X _25402_/S vssd1 vssd1 vccd1 vccd1 _25395_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27133_ _27133_/CLK _27133_/D vssd1 vssd1 vccd1 vccd1 _27133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24345_ _24345_/A vssd1 vssd1 vccd1 vccd1 _27455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21557_ _21545_/X _21546_/X _21547_/X _21548_/X _21549_/X _21550_/X vssd1 vssd1 vccd1
+ vccd1 _21558_/A sky130_fd_sc_hd__mux4_1
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20508_ _20496_/X _20497_/X _20498_/X _20499_/X _20500_/X _20501_/X vssd1 vssd1 vccd1
+ vccd1 _20509_/A sky130_fd_sc_hd__mux4_1
X_27064_ _23024_/X _27064_/D vssd1 vssd1 vccd1 vccd1 _27064_/Q sky130_fd_sc_hd__dfxtp_1
X_24276_ _16221_/X _16223_/Y _16224_/X _24273_/X vssd1 vssd1 vccd1 vccd1 _27413_/D
+ sky130_fd_sc_hd__o31a_1
X_21488_ _21488_/A vssd1 vssd1 vccd1 vccd1 _21488_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26015_ _27416_/CLK _26015_/D vssd1 vssd1 vccd1 vccd1 _26015_/Q sky130_fd_sc_hd__dfxtp_1
X_23227_ _23227_/A vssd1 vssd1 vccd1 vccd1 _27149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20439_ _20439_/A vssd1 vssd1 vccd1 vccd1 _20439_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23158_ _23158_/A vssd1 vssd1 vccd1 vccd1 _27118_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22109_ _22175_/A vssd1 vssd1 vccd1 vccd1 _22109_/X sky130_fd_sc_hd__clkbuf_1
X_15980_ _15980_/A vssd1 vssd1 vccd1 vccd1 _15985_/A sky130_fd_sc_hd__buf_6
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23089_ _23089_/A vssd1 vssd1 vccd1 vccd1 _27088_/D sky130_fd_sc_hd__clkbuf_1
X_27966_ _27966_/A _15865_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
XFILLER_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14931_ _14942_/A vssd1 vssd1 vccd1 vccd1 _14940_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_88_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26917_ _22514_/X _26917_/D vssd1 vssd1 vccd1 vccd1 _26917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17650_ _17492_/X _25896_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _17651_/A sky130_fd_sc_hd__mux2_1
X_14862_ _26500_/Q _13389_/X _14868_/S vssd1 vssd1 vccd1 vccd1 _14863_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26848_ _22276_/X _26848_/D vssd1 vssd1 vccd1 vccd1 _26848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13813_ _26856_/Q _13806_/X _13807_/X _13812_/Y vssd1 vssd1 vccd1 vccd1 _26856_/D
+ sky130_fd_sc_hd__a31o_1
X_16601_ _16309_/Y _16902_/A _16600_/Y _16309_/A vssd1 vssd1 vccd1 vccd1 _16604_/A
+ sky130_fd_sc_hd__o31a_1
X_17581_ _17581_/A vssd1 vssd1 vccd1 vccd1 _25865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26779_ _22034_/X _26779_/D vssd1 vssd1 vccd1 vccd1 _26779_/Q sky130_fd_sc_hd__dfxtp_1
X_14793_ _14791_/X _26528_/Q _14805_/S vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19320_ _26958_/Q _26926_/Q _26894_/Q _26862_/Q _19208_/X _19253_/X vssd1 vssd1 vccd1
+ vccd1 _19320_/X sky130_fd_sc_hd__mux4_1
X_16532_ _16845_/A _16623_/B vssd1 vssd1 vccd1 vccd1 _16534_/A sky130_fd_sc_hd__nand2_1
X_13744_ _26881_/Q _13737_/X _13732_/X _13743_/Y vssd1 vssd1 vccd1 vccd1 _26881_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19251_ _26699_/Q _26667_/Q _26635_/Q _26603_/Q _19179_/X _19227_/X vssd1 vssd1 vccd1
+ vccd1 _19251_/X sky130_fd_sc_hd__mux4_2
X_16463_ _16470_/A _16471_/B vssd1 vssd1 vccd1 vccd1 _16692_/C sky130_fd_sc_hd__xnor2_1
X_13675_ _13691_/A vssd1 vssd1 vccd1 vccd1 _13759_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18202_ _18202_/A _18156_/X vssd1 vssd1 vccd1 vccd1 _18202_/X sky130_fd_sc_hd__or2b_1
X_15414_ _26263_/Q _13328_/X _15418_/S vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__mux2_1
X_19182_ _26952_/Q _26920_/Q _26888_/Q _26856_/Q _19044_/X _19116_/X vssd1 vssd1 vccd1
+ vccd1 _19182_/X sky130_fd_sc_hd__mux4_2
XFILLER_188_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16394_ _16745_/B _16396_/B vssd1 vssd1 vccd1 vccd1 _16394_/X sky130_fd_sc_hd__or2_1
X_18133_ _26693_/Q _26661_/Q _26629_/Q _26597_/Q _18036_/X _18106_/X vssd1 vssd1 vccd1
+ vccd1 _18134_/A sky130_fd_sc_hd__mux4_2
XFILLER_106_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15345_ _15345_/A vssd1 vssd1 vccd1 vccd1 _26294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18064_ _17972_/X _18056_/X _18063_/X _17932_/X vssd1 vssd1 vccd1 vccd1 _18077_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ _26324_/Q _13337_/X _15284_/S vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17015_ _17291_/A vssd1 vssd1 vccd1 vccd1 _17015_/X sky130_fd_sc_hd__clkbuf_4
X_14227_ _26718_/Q _14225_/X _14220_/X _14226_/Y vssd1 vssd1 vccd1 vccd1 _26718_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14158_ _14335_/A _14158_/B vssd1 vssd1 vccd1 vccd1 _14158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _27293_/Q _13109_/B vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__and2_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _26769_/Q _14076_/X _14080_/X _14088_/Y vssd1 vssd1 vccd1 vccd1 _26769_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _18966_/A vssd1 vssd1 vccd1 vccd1 _26046_/D sky130_fd_sc_hd__clkbuf_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _17897_/X _17907_/X _17911_/X _17916_/X _17856_/X vssd1 vssd1 vccd1 vccd1
+ _17918_/C sky130_fd_sc_hd__a221o_1
XFILLER_117_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18897_ _18897_/A vssd1 vssd1 vccd1 vccd1 _19445_/A sky130_fd_sc_hd__buf_4
XFILLER_152_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17848_ _18418_/A vssd1 vssd1 vccd1 vccd1 _17848_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_187_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17779_ _18150_/A vssd1 vssd1 vccd1 vccd1 _17779_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19518_ _19431_/X _19517_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _19518_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20790_ _21143_/A vssd1 vssd1 vccd1 vccd1 _20864_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19449_ _19440_/X _19443_/X _19447_/X _19448_/X _19360_/X vssd1 vssd1 vccd1 vccd1
+ _19450_/C sky130_fd_sc_hd__a221o_1
XFILLER_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22460_ _22508_/A vssd1 vssd1 vccd1 vccd1 _22460_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21411_ _21583_/A vssd1 vssd1 vccd1 vccd1 _21477_/A sky130_fd_sc_hd__clkbuf_2
X_22391_ _22385_/X _22386_/X _22387_/X _22388_/X _22389_/X _22390_/X vssd1 vssd1 vccd1
+ vccd1 _22392_/A sky130_fd_sc_hd__mux4_1
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24130_ _24186_/A vssd1 vssd1 vccd1 vccd1 _24175_/A sky130_fd_sc_hd__clkbuf_2
X_21342_ _21390_/A vssd1 vssd1 vccd1 vccd1 _21342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24061_ _24061_/A _24061_/B vssd1 vssd1 vccd1 vccd1 _24062_/A sky130_fd_sc_hd__and2_1
XFILLER_200_1073 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21273_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21273_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23012_ _25638_/A vssd1 vssd1 vccd1 vccd1 _23012_/X sky130_fd_sc_hd__clkbuf_1
X_20224_ _20216_/X _20217_/X _20218_/X _20219_/X _20220_/X _20221_/X vssd1 vssd1 vccd1
+ vccd1 _20225_/A sky130_fd_sc_hd__mux4_1
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27820_ _25718_/X _27820_/D vssd1 vssd1 vccd1 vccd1 _27820_/Q sky130_fd_sc_hd__dfxtp_1
X_20155_ _20155_/A vssd1 vssd1 vccd1 vccd1 _20155_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27751_ _27751_/CLK _27751_/D vssd1 vssd1 vccd1 vccd1 _27751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20086_ _20076_/X _20077_/X _20078_/X _20079_/X _20081_/X _20083_/X vssd1 vssd1 vccd1
+ vccd1 _20087_/A sky130_fd_sc_hd__mux4_1
X_24963_ _27669_/Q _24838_/A _24962_/Y _24663_/A vssd1 vssd1 vccd1 vccd1 _27669_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26702_ _21772_/X _26702_/D vssd1 vssd1 vccd1 vccd1 _26702_/Q sky130_fd_sc_hd__dfxtp_1
X_23914_ _25928_/Q _25994_/Q _25827_/Q _26026_/Q _23899_/X _23882_/X vssd1 vssd1 vccd1
+ vccd1 _23914_/X sky130_fd_sc_hd__mux4_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27682_ _27682_/CLK _27682_/D vssd1 vssd1 vccd1 vccd1 _27973_/A sky130_fd_sc_hd__dfxtp_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24894_ _24913_/A _24894_/B vssd1 vssd1 vccd1 vccd1 _24894_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26633_ _21526_/X _26633_/D vssd1 vssd1 vccd1 vccd1 _26633_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23845_ _27075_/Q _27107_/Q _23845_/S vssd1 vssd1 vccd1 vccd1 _23845_/X sky130_fd_sc_hd__mux2_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26564_ _21284_/X _26564_/D vssd1 vssd1 vccd1 vccd1 _26564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23776_ _23740_/X _23774_/X _23775_/X _23768_/X vssd1 vssd1 vccd1 vccd1 _27272_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20988_ _20988_/A vssd1 vssd1 vccd1 vccd1 _20988_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25515_ _24767_/A _25504_/X _25511_/Y _25514_/X _25497_/X vssd1 vssd1 vccd1 vccd1
+ _27766_/D sky130_fd_sc_hd__a221oi_1
XFILLER_198_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22727_ _22716_/X _22718_/X _22720_/X _22722_/X _22723_/X _22724_/X vssd1 vssd1 vccd1
+ vccd1 _22728_/A sky130_fd_sc_hd__mux4_1
XFILLER_201_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26495_ _21048_/X _26495_/D vssd1 vssd1 vccd1 vccd1 _26495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13460_ _13874_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13460_/Y sky130_fd_sc_hd__nor2_1
X_25446_ _25466_/A vssd1 vssd1 vccd1 vccd1 _25446_/X sky130_fd_sc_hd__clkbuf_2
X_22658_ _22658_/A vssd1 vssd1 vccd1 vccd1 _22658_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21609_ _21599_/X _21600_/X _21601_/X _21602_/X _21603_/X _21604_/X vssd1 vssd1 vccd1
+ vccd1 _21610_/A sky130_fd_sc_hd__mux4_1
XFILLER_127_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25377_ _25377_/A vssd1 vssd1 vccd1 vccd1 _27728_/D sky130_fd_sc_hd__clkbuf_1
X_13391_ _13391_/A vssd1 vssd1 vccd1 vccd1 _26980_/D sky130_fd_sc_hd__clkbuf_1
X_22589_ _22577_/X _22578_/X _22579_/X _22580_/X _22581_/X _22582_/X vssd1 vssd1 vccd1
+ vccd1 _22590_/A sky130_fd_sc_hd__mux4_1
XFILLER_154_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27116_ _27214_/CLK _27116_/D vssd1 vssd1 vccd1 vccd1 _27116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ _15130_/A vssd1 vssd1 vccd1 vccd1 _26389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_782 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_601 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24328_ _27548_/Q _24328_/B vssd1 vssd1 vccd1 vccd1 _24329_/A sky130_fd_sc_hd__and2_1
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27047_ _22968_/X _27047_/D vssd1 vssd1 vccd1 vccd1 _27047_/Q sky130_fd_sc_hd__dfxtp_1
X_15061_ _15061_/A vssd1 vssd1 vccd1 vccd1 _26420_/D sky130_fd_sc_hd__clkbuf_1
X_24259_ _24259_/A _24287_/B vssd1 vssd1 vccd1 vccd1 _24260_/A sky130_fd_sc_hd__and2_1
X_14012_ _16243_/A vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18820_ _27601_/Q vssd1 vssd1 vccd1 vccd1 _19387_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_862 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18751_ _26036_/Q _17760_/X _18757_/S vssd1 vssd1 vccd1 vccd1 _18752_/A sky130_fd_sc_hd__mux2_1
X_15963_ _15967_/A vssd1 vssd1 vccd1 vccd1 _15963_/Y sky130_fd_sc_hd__inv_2
X_27949_ _27949_/A _15927_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17702_ _27416_/Q vssd1 vssd1 vccd1 vccd1 _17702_/X sky130_fd_sc_hd__clkbuf_2
X_14914_ _14750_/X _26477_/Q _14918_/S vssd1 vssd1 vccd1 vccd1 _14915_/A sky130_fd_sc_hd__mux2_1
X_18682_ _18682_/A vssd1 vssd1 vccd1 vccd1 _26005_/D sky130_fd_sc_hd__clkbuf_1
X_15894_ _15894_/A vssd1 vssd1 vccd1 vccd1 _15899_/A sky130_fd_sc_hd__buf_4
X_17633_ _17633_/A vssd1 vssd1 vccd1 vccd1 _25888_/D sky130_fd_sc_hd__clkbuf_1
X_14845_ _14845_/A vssd1 vssd1 vccd1 vccd1 _26508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17564_ _17586_/A vssd1 vssd1 vccd1 vccd1 _17573_/S sky130_fd_sc_hd__clkbuf_2
X_14776_ _14792_/A vssd1 vssd1 vccd1 vccd1 _14789_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19303_ _26157_/Q _26093_/Q _27021_/Q _26989_/Q _18923_/A _18926_/A vssd1 vssd1 vccd1
+ vccd1 _19304_/B sky130_fd_sc_hd__mux4_2
X_13727_ _13740_/A vssd1 vssd1 vccd1 vccd1 _13738_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16515_ _27398_/Q _16094_/A _16314_/X _14740_/A vssd1 vssd1 vccd1 vccd1 _16515_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17495_ _27430_/Q vssd1 vssd1 vccd1 vccd1 _17495_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19234_ _19231_/X _19232_/X _19346_/S vssd1 vssd1 vccd1 vccd1 _19234_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13658_ _26912_/Q _13653_/X _13656_/X _13657_/Y vssd1 vssd1 vccd1 vccd1 _26912_/D
+ sky130_fd_sc_hd__a31o_1
X_16446_ _16036_/X _16162_/Y _16445_/X _16164_/X vssd1 vssd1 vccd1 vccd1 _16446_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_108_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19165_ _19165_/A vssd1 vssd1 vccd1 vccd1 _19165_/X sky130_fd_sc_hd__buf_2
X_16377_ _16749_/B vssd1 vssd1 vccd1 vccd1 _16751_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13589_ _13857_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15328_ _26300_/Q _13414_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15329_/A sky130_fd_sc_hd__mux2_1
X_18116_ _18020_/X _18115_/X _18070_/X vssd1 vssd1 vccd1 vccd1 _18116_/X sky130_fd_sc_hd__o21a_1
XFILLER_173_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19096_ _26148_/Q _26084_/Q _27012_/Q _26980_/Q _19049_/X _19070_/X vssd1 vssd1 vccd1
+ vccd1 _19097_/B sky130_fd_sc_hd__mux4_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18047_ _26529_/Q _26497_/Q _26465_/Q _27041_/Q _17964_/X _17986_/X vssd1 vssd1 vccd1
+ vccd1 _18047_/X sky130_fd_sc_hd__mux4_1
X_15259_ _15259_/A vssd1 vssd1 vccd1 vccd1 _26331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19998_ _19988_/X _19989_/X _19990_/X _19991_/X _19994_/X _19997_/X vssd1 vssd1 vccd1
+ vccd1 _19999_/A sky130_fd_sc_hd__mux4_1
XFILLER_115_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18949_ _19208_/A vssd1 vssd1 vccd1 vccd1 _19482_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21960_ _21960_/A vssd1 vssd1 vccd1 vccd1 _21960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20911_ _20905_/X _20906_/X _20907_/X _20908_/X _20909_/X _20910_/X vssd1 vssd1 vccd1
+ vccd1 _20912_/A sky130_fd_sc_hd__mux4_1
X_21891_ _21879_/X _21880_/X _21881_/X _21882_/X _21883_/X _21884_/X vssd1 vssd1 vccd1
+ vccd1 _21892_/A sky130_fd_sc_hd__mux4_1
XFILLER_199_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23630_ _27229_/Q vssd1 vssd1 vccd1 vccd1 _25018_/A sky130_fd_sc_hd__buf_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20842_ _20832_/X _20833_/X _20834_/X _20835_/X _20836_/X _20837_/X vssd1 vssd1 vccd1
+ vccd1 _20843_/A sky130_fd_sc_hd__mux4_1
XFILLER_74_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23561_ _23561_/A vssd1 vssd1 vccd1 vccd1 _27209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20773_ _20773_/A vssd1 vssd1 vccd1 vccd1 _20773_/X sky130_fd_sc_hd__clkbuf_1
X_25300_ _27510_/Q _27509_/Q _27508_/Q _27507_/Q _25310_/A vssd1 vssd1 vccd1 vccd1
+ _25300_/X sky130_fd_sc_hd__o41a_1
XFILLER_167_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22512_ _22512_/A vssd1 vssd1 vccd1 vccd1 _22512_/X sky130_fd_sc_hd__clkbuf_1
X_26280_ _20293_/X _26280_/D vssd1 vssd1 vccd1 vccd1 _26280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23492_ input28/X _23482_/X _23491_/X _23487_/X vssd1 vssd1 vccd1 vccd1 _27189_/D
+ sky130_fd_sc_hd__o211a_1
X_25231_ _27704_/Q _25223_/X _25230_/Y _25214_/X vssd1 vssd1 vccd1 vccd1 _27704_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22443_ _22433_/X _22434_/X _22435_/X _22436_/X _22438_/X _22440_/X vssd1 vssd1 vccd1
+ vccd1 _22444_/A sky130_fd_sc_hd__mux4_1
XFILLER_129_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25162_ _25162_/A _25162_/B vssd1 vssd1 vccd1 vccd1 _25165_/A sky130_fd_sc_hd__nand2_1
XFILLER_175_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22374_ _22422_/A vssd1 vssd1 vccd1 vccd1 _22374_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24113_ _27404_/Q _24117_/B vssd1 vssd1 vccd1 vccd1 _24114_/A sky130_fd_sc_hd__and2_1
X_21325_ _21583_/A vssd1 vssd1 vccd1 vccd1 _21391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25093_ _25926_/Q _25992_/Q _25825_/Q _26024_/Q _25018_/A _25070_/X vssd1 vssd1 vccd1
+ vccd1 _25093_/X sky130_fd_sc_hd__mux4_1
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24044_ _25943_/Q _26009_/Q _25842_/Q _26041_/Q _23777_/A _23744_/A vssd1 vssd1 vccd1
+ vccd1 _24044_/X sky130_fd_sc_hd__mux4_1
X_21256_ _21304_/A vssd1 vssd1 vccd1 vccd1 _21256_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20207_ _20207_/A vssd1 vssd1 vccd1 vccd1 _20207_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21187_ _21179_/X _21180_/X _21181_/X _21182_/X _21183_/X _21184_/X vssd1 vssd1 vccd1
+ vccd1 _21188_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_28016__482 vssd1 vssd1 vccd1 vccd1 _28016__482/HI _28016_/A sky130_fd_sc_hd__conb_1
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27803_ _25666_/X _27803_/D vssd1 vssd1 vccd1 vccd1 _27803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20138_ _20130_/X _20131_/X _20132_/X _20133_/X _20134_/X _20135_/X vssd1 vssd1 vccd1
+ vccd1 _20139_/A sky130_fd_sc_hd__mux4_1
X_25995_ _25995_/CLK _25995_/D vssd1 vssd1 vccd1 vccd1 _25995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12960_/A vssd1 vssd1 vccd1 vccd1 _27817_/D sky130_fd_sc_hd__clkbuf_1
X_27734_ _27735_/CLK _27734_/D vssd1 vssd1 vccd1 vccd1 _27734_/Q sky130_fd_sc_hd__dfxtp_1
X_20069_ _20069_/A vssd1 vssd1 vccd1 vccd1 _20069_/X sky130_fd_sc_hd__clkbuf_1
X_24946_ _24947_/A _24947_/B vssd1 vssd1 vccd1 vccd1 _24954_/C sky130_fd_sc_hd__and2_1
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_482 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24877_ _24877_/A _24880_/C vssd1 vssd1 vccd1 vccd1 _24878_/B sky130_fd_sc_hd__xnor2_1
X_27665_ _27668_/CLK _27665_/D vssd1 vssd1 vccd1 vccd1 _27665_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 _20695_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 _18196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14671_/A vssd1 vssd1 vccd1 vccd1 _14630_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _19161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26616_ _21468_/X _26616_/D vssd1 vssd1 vccd1 vccd1 _26616_/Q sky130_fd_sc_hd__dfxtp_1
X_23828_ _25919_/Q _25985_/Q _25818_/Q _26017_/Q _23804_/X _23786_/X vssd1 vssd1 vccd1
+ vccd1 _23828_/X sky130_fd_sc_hd__mux4_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27596_ _27597_/CLK _27596_/D vssd1 vssd1 vccd1 vccd1 _27596_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_334 _13122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _13414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_356 _14718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _26817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14561_ _15723_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14561_/Y sky130_fd_sc_hd__nor2_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26547_ _21224_/X _26547_/D vssd1 vssd1 vccd1 vccd1 _26547_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_378 _24386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23759_ _23753_/X _23756_/X _23797_/S vssd1 vssd1 vccd1 vccd1 _23759_/X sky130_fd_sc_hd__mux2_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _16451_/A vssd1 vssd1 vccd1 vccd1 _13902_/A sky130_fd_sc_hd__clkbuf_2
X_16300_ _16583_/A _16648_/B vssd1 vssd1 vccd1 vccd1 _16301_/D sky130_fd_sc_hd__nand2_1
XFILLER_41_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _25833_/Q _26032_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17280_/X sky130_fd_sc_hd__mux2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14510_/A vssd1 vssd1 vccd1 vccd1 _14492_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26478_ _20988_/X _26478_/D vssd1 vssd1 vccd1 vccd1 _26478_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _27527_/Q _15992_/A vssd1 vssd1 vccd1 vccd1 _16231_/X sky130_fd_sc_hd__or2b_1
X_13443_ _26967_/Q _13435_/X _13429_/X _13442_/Y vssd1 vssd1 vccd1 vccd1 _26967_/D
+ sky130_fd_sc_hd__a31o_1
X_25429_ _25429_/A vssd1 vssd1 vccd1 vccd1 _27752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16162_ _16420_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16162_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13374_ _26985_/Q _13373_/X _13383_/S vssd1 vssd1 vccd1 vccd1 _13375_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15113_ _15113_/A vssd1 vssd1 vccd1 vccd1 _26396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16093_ _16619_/A vssd1 vssd1 vccd1 vccd1 _16093_/X sky130_fd_sc_hd__buf_2
XFILLER_155_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15044_ _26426_/Q _15040_/X _14966_/B _15043_/Y vssd1 vssd1 vccd1 vccd1 _26426_/D
+ sky130_fd_sc_hd__a31o_1
X_19921_ _19989_/A vssd1 vssd1 vccd1 vccd1 _19921_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19852_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19852_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _18772_/X _18786_/X _18799_/X _18801_/X _24407_/A vssd1 vssd1 vccd1 vccd1
+ _18842_/B sky130_fd_sc_hd__a221o_1
XFILLER_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19783_ _19815_/A vssd1 vssd1 vccd1 vccd1 _19783_/X sky130_fd_sc_hd__clkbuf_1
X_16995_ _25912_/Q _25978_/Q _17382_/S vssd1 vssd1 vccd1 vccd1 _16996_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18734_ _18734_/A vssd1 vssd1 vccd1 vccd1 _26028_/D sky130_fd_sc_hd__clkbuf_1
X_15946_ _15949_/A vssd1 vssd1 vccd1 vccd1 _15946_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18665_ _18676_/A vssd1 vssd1 vccd1 vccd1 _18674_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _15881_/A vssd1 vssd1 vccd1 vccd1 _15877_/Y sky130_fd_sc_hd__inv_2
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17616_ _17616_/A vssd1 vssd1 vccd1 vccd1 _25880_/D sky130_fd_sc_hd__clkbuf_1
X_14828_ _14828_/A vssd1 vssd1 vccd1 vccd1 _26516_/D sky130_fd_sc_hd__clkbuf_1
X_18596_ _27540_/Q _27519_/Q vssd1 vssd1 vccd1 vccd1 _18613_/A sky130_fd_sc_hd__nand2_1
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17547_ _17447_/X _25850_/Q _17551_/S vssd1 vssd1 vccd1 vccd1 _17548_/A sky130_fd_sc_hd__mux2_1
X_14759_ _14759_/A vssd1 vssd1 vccd1 vccd1 _14759_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17478_ _17478_/A vssd1 vssd1 vccd1 vccd1 _25827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19217_ _19555_/A _19217_/B vssd1 vssd1 vccd1 vccd1 _19217_/X sky130_fd_sc_hd__or2_1
X_16429_ _16359_/A _16447_/C _16447_/D _16369_/X vssd1 vssd1 vccd1 vccd1 _16430_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_146_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19148_ _19287_/A vssd1 vssd1 vccd1 vccd1 _19148_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19079_ _26531_/Q _26499_/Q _26467_/Q _27043_/Q _18984_/X _19032_/X vssd1 vssd1 vccd1
+ vccd1 _19079_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_402 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21110_ _21126_/A vssd1 vssd1 vccd1 vccd1 _21110_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22090_ _22162_/A vssd1 vssd1 vccd1 vccd1 _22090_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21041_ _21041_/A vssd1 vssd1 vccd1 vccd1 _21041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24800_ _24800_/A _24800_/B vssd1 vssd1 vccd1 vccd1 _24800_/Y sky130_fd_sc_hd__nand2_1
X_25780_ _25780_/A vssd1 vssd1 vccd1 vccd1 _27845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22992_ _22992_/A vssd1 vssd1 vccd1 vccd1 _22992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24731_ _27193_/Q _25474_/A vssd1 vssd1 vccd1 vccd1 _24731_/X sky130_fd_sc_hd__or2_1
X_21943_ _21930_/X _21932_/X _21934_/X _21936_/X _21937_/X _21938_/X vssd1 vssd1 vccd1
+ vccd1 _21944_/A sky130_fd_sc_hd__mux4_1
X_27450_ _27450_/CLK _27450_/D vssd1 vssd1 vccd1 vccd1 _27450_/Q sky130_fd_sc_hd__dfxtp_1
X_24662_ _27167_/Q _24671_/B vssd1 vssd1 vccd1 vccd1 _24662_/X sky130_fd_sc_hd__or2_1
X_21874_ _21874_/A vssd1 vssd1 vccd1 vccd1 _21874_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26401_ _20715_/X _26401_/D vssd1 vssd1 vccd1 vccd1 _26401_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23613_ _23617_/A _23613_/B vssd1 vssd1 vccd1 vccd1 _23614_/A sky130_fd_sc_hd__and2_1
X_20825_ _20825_/A vssd1 vssd1 vccd1 vccd1 _20825_/X sky130_fd_sc_hd__clkbuf_1
X_27381_ _27383_/CLK _27381_/D vssd1 vssd1 vccd1 vccd1 _27381_/Q sky130_fd_sc_hd__dfxtp_1
X_24593_ _24593_/A vssd1 vssd1 vccd1 vccd1 _27556_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26332_ _20475_/X _26332_/D vssd1 vssd1 vccd1 vccd1 _26332_/Q sky130_fd_sc_hd__dfxtp_1
X_23544_ _23544_/A vssd1 vssd1 vccd1 vccd1 _27204_/D sky130_fd_sc_hd__clkbuf_1
X_20756_ _20772_/A vssd1 vssd1 vccd1 vccd1 _20756_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26263_ _20229_/X _26263_/D vssd1 vssd1 vccd1 vccd1 _26263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23475_ input21/X _23469_/X _23473_/X _23474_/X vssd1 vssd1 vccd1 vccd1 _27182_/D
+ sky130_fd_sc_hd__o211a_1
X_20687_ _20687_/A vssd1 vssd1 vccd1 vccd1 _20687_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25214_ _25297_/A vssd1 vssd1 vccd1 vccd1 _25214_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_28002_ _28002_/A _15878_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_22426_ _22426_/A vssd1 vssd1 vccd1 vccd1 _22426_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26194_ _19987_/X _26194_/D vssd1 vssd1 vccd1 vccd1 _26194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25145_ _27524_/Q _27492_/Q vssd1 vssd1 vccd1 vccd1 _25147_/A sky130_fd_sc_hd__and2_1
X_22357_ _22347_/X _22348_/X _22349_/X _22350_/X _22352_/X _22354_/X vssd1 vssd1 vccd1
+ vccd1 _22358_/A sky130_fd_sc_hd__mux4_1
XFILLER_156_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21308_ _22616_/A vssd1 vssd1 vccd1 vccd1 _21653_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25076_ _27974_/A _25074_/X _25104_/S vssd1 vssd1 vccd1 vccd1 _25077_/A sky130_fd_sc_hd__mux2_1
X_13090_ _13529_/A vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__clkbuf_2
X_22288_ _22336_/A vssd1 vssd1 vccd1 vccd1 _22288_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24027_ _27094_/Q _24001_/X _24002_/X _27126_/Q _24003_/X vssd1 vssd1 vccd1 vccd1
+ _24027_/X sky130_fd_sc_hd__a221o_1
X_21239_ _21585_/A vssd1 vssd1 vccd1 vccd1 _21304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _15800_/A vssd1 vssd1 vccd1 vccd1 _26099_/D sky130_fd_sc_hd__clkbuf_1
X_13992_ _14363_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16780_ _16780_/A _16780_/B _16767_/A vssd1 vssd1 vccd1 vccd1 _16780_/X sky130_fd_sc_hd__or3b_1
X_25978_ _27076_/CLK _25978_/D vssd1 vssd1 vccd1 vccd1 _25978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _26126_/Q _15721_/X _15727_/X _15730_/Y vssd1 vssd1 vccd1 vccd1 _26126_/D
+ sky130_fd_sc_hd__a31o_1
X_12943_ _23598_/A vssd1 vssd1 vccd1 vccd1 _12952_/B sky130_fd_sc_hd__clkbuf_1
X_27717_ _27772_/CLK _27717_/D vssd1 vssd1 vccd1 vccd1 _27717_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24929_ _27662_/Q _24909_/X _24928_/Y _24914_/X vssd1 vssd1 vccd1 vccd1 _27662_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18450_ _26707_/Q _26675_/Q _26643_/Q _26611_/Q _17782_/X _18005_/X vssd1 vssd1 vccd1
+ vccd1 _18451_/A sky130_fd_sc_hd__mux4_2
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _22546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27648_ _27667_/CLK _27648_/D vssd1 vssd1 vccd1 vccd1 _27648_/Q sky130_fd_sc_hd__dfxtp_1
X_15662_ _15662_/A vssd1 vssd1 vccd1 vccd1 _26153_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _23991_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ input4/X vssd1 vssd1 vccd1 vccd1 _25639_/A sky130_fd_sc_hd__buf_4
XANTENNA_142 _13038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14613_ _26589_/Q _14602_/X _14605_/X _14612_/Y vssd1 vssd1 vccd1 vccd1 _26589_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA_153 _13319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18381_ _26832_/Q _26800_/Q _26768_/Q _26736_/Q _18358_/X _18380_/X vssd1 vssd1 vccd1
+ vccd1 _18381_/X sky130_fd_sc_hd__mux4_1
X_15593_ _26183_/Q _14769_/A _15595_/S vssd1 vssd1 vccd1 vccd1 _15594_/A sky130_fd_sc_hd__mux2_1
XANTENNA_164 _13389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _14448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27579_ _27584_/CLK _27579_/D vssd1 vssd1 vccd1 vccd1 _27579_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _14471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17332_ _17299_/X _17326_/X _17329_/X _17331_/X vssd1 vssd1 vccd1 vccd1 _17332_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_197 _14493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14544_ _14552_/A vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14475_ _16495_/A vssd1 vssd1 vccd1 vccd1 _15741_/A sky130_fd_sc_hd__buf_2
X_17263_ _17263_/A vssd1 vssd1 vccd1 vccd1 _27936_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ _18995_/X _18998_/X _19001_/X _18854_/X _18880_/X vssd1 vssd1 vccd1 vccd1
+ _19011_/B sky130_fd_sc_hd__a221o_2
X_13426_ _15623_/B vssd1 vssd1 vccd1 vccd1 _15335_/A sky130_fd_sc_hd__buf_4
X_16214_ _16180_/X _16209_/X _16211_/Y _16212_/X _16213_/X vssd1 vssd1 vccd1 vccd1
+ _16388_/A sky130_fd_sc_hd__o41a_1
X_17194_ _17155_/X _17194_/B vssd1 vssd1 vccd1 vccd1 _17194_/X sky130_fd_sc_hd__and2b_1
X_16145_ _16143_/Y _16119_/X _16121_/X _16563_/A _16144_/Y vssd1 vssd1 vccd1 vccd1
+ _24302_/A sky130_fd_sc_hd__o221a_1
X_13357_ _14747_/A vssd1 vssd1 vccd1 vccd1 _13357_/X sky130_fd_sc_hd__buf_2
XFILLER_6_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16076_ _16076_/A vssd1 vssd1 vccd1 vccd1 _16077_/A sky130_fd_sc_hd__clkbuf_2
X_13288_ _13288_/A vssd1 vssd1 vccd1 vccd1 _27016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15027_ _26433_/Q _15015_/X _15016_/X _15026_/Y vssd1 vssd1 vccd1 vccd1 _26433_/D
+ sky130_fd_sc_hd__a31o_1
X_19904_ _25726_/A vssd1 vssd1 vccd1 vccd1 _19977_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19835_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19835_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19766_ _19814_/A vssd1 vssd1 vccd1 vccd1 _19766_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16978_ _24435_/A vssd1 vssd1 vccd1 vccd1 _24624_/B sky130_fd_sc_hd__buf_2
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_18717_ _18717_/A vssd1 vssd1 vccd1 vccd1 _26020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15929_ _15930_/A vssd1 vssd1 vccd1 vccd1 _15929_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19697_ _19729_/A vssd1 vssd1 vccd1 vccd1 _19697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18648_ _25990_/Q _17715_/X _18652_/S vssd1 vssd1 vccd1 vccd1 _18649_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18579_ _26425_/Q _26393_/Q _26361_/Q _26329_/Q _17996_/X _18486_/X vssd1 vssd1 vccd1
+ vccd1 _18579_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20610_ _20598_/X _20599_/X _20600_/X _20601_/X _20603_/X _20605_/X vssd1 vssd1 vccd1
+ vccd1 _20611_/A sky130_fd_sc_hd__mux4_1
X_21590_ _21590_/A vssd1 vssd1 vccd1 vccd1 _21590_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20541_ _20541_/A vssd1 vssd1 vccd1 vccd1 _20541_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23260_ _27729_/Q vssd1 vssd1 vccd1 vccd1 _23260_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20472_ _20464_/X _20465_/X _20466_/X _20467_/X _20468_/X _20469_/X vssd1 vssd1 vccd1
+ vccd1 _20473_/A sky130_fd_sc_hd__mux4_1
X_22211_ _22194_/X _22196_/X _22198_/X _22200_/X _22201_/X _22202_/X vssd1 vssd1 vccd1
+ vccd1 _22212_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23191_ _17434_/X _27133_/Q _23193_/S vssd1 vssd1 vccd1 vccd1 _23192_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22142_ _22174_/A vssd1 vssd1 vccd1 vccd1 _22142_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22073_ _22067_/X _22068_/X _22069_/X _22070_/X _22071_/X _22072_/X vssd1 vssd1 vccd1
+ vccd1 _22074_/A sky130_fd_sc_hd__mux4_1
X_26950_ _22640_/X _26950_/D vssd1 vssd1 vccd1 vccd1 _26950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25901_ _25901_/CLK _25901_/D vssd1 vssd1 vccd1 vccd1 _25901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21024_ _21040_/A vssd1 vssd1 vccd1 vccd1 _21024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26881_ _22394_/X _26881_/D vssd1 vssd1 vccd1 vccd1 _26881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25832_ _27088_/CLK _25832_/D vssd1 vssd1 vccd1 vccd1 _25832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25763_ _25763_/A vssd1 vssd1 vccd1 vccd1 _27837_/D sky130_fd_sc_hd__clkbuf_1
X_22975_ _25655_/A vssd1 vssd1 vccd1 vccd1 _25636_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27502_ _27623_/CLK _27502_/D vssd1 vssd1 vccd1 vccd1 _27502_/Q sky130_fd_sc_hd__dfxtp_1
X_21926_ _21926_/A vssd1 vssd1 vccd1 vccd1 _21926_/X sky130_fd_sc_hd__clkbuf_1
X_24714_ _24771_/A vssd1 vssd1 vccd1 vccd1 _24714_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25694_ _25710_/A vssd1 vssd1 vccd1 vccd1 _25694_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27433_ _27435_/CLK _27433_/D vssd1 vssd1 vccd1 vccd1 _27433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24645_ _25540_/A vssd1 vssd1 vccd1 vccd1 _24658_/B sky130_fd_sc_hd__clkbuf_1
X_21857_ _21844_/X _21846_/X _21848_/X _21850_/X _21851_/X _21852_/X vssd1 vssd1 vccd1
+ vccd1 _21858_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _20791_/X _20795_/X _20799_/X _20803_/X _20804_/X _20805_/X vssd1 vssd1 vccd1
+ vccd1 _20809_/A sky130_fd_sc_hd__mux4_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24576_ _27649_/Q _24576_/B vssd1 vssd1 vccd1 vccd1 _24577_/A sky130_fd_sc_hd__and2_1
X_27364_ _27365_/CLK _27364_/D vssd1 vssd1 vccd1 vccd1 _27364_/Q sky130_fd_sc_hd__dfxtp_1
X_21788_ _21788_/A vssd1 vssd1 vccd1 vccd1 _21788_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26315_ _20415_/X _26315_/D vssd1 vssd1 vccd1 vccd1 _26315_/Q sky130_fd_sc_hd__dfxtp_1
X_23527_ _23527_/A vssd1 vssd1 vccd1 vccd1 _27199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27295_ _27295_/CLK _27295_/D vssd1 vssd1 vccd1 vccd1 _27295_/Q sky130_fd_sc_hd__dfxtp_1
X_20739_ _20771_/A vssd1 vssd1 vccd1 vccd1 _20739_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14260_ _26708_/Q _14256_/X _14258_/X _14259_/Y vssd1 vssd1 vccd1 vccd1 _26708_/D
+ sky130_fd_sc_hd__a31o_1
X_26246_ _20173_/X _26246_/D vssd1 vssd1 vccd1 vccd1 _26246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23458_ _23485_/A vssd1 vssd1 vccd1 vccd1 _23470_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13211_ _27039_/Q _13210_/X _13229_/S vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__mux2_1
X_22409_ _22401_/X _22402_/X _22403_/X _22404_/X _22405_/X _22406_/X vssd1 vssd1 vccd1
+ vccd1 _22410_/A sky130_fd_sc_hd__mux4_1
X_14191_ _26732_/Q _14186_/X _14181_/X _14190_/Y vssd1 vssd1 vccd1 vccd1 _26732_/D
+ sky130_fd_sc_hd__a31o_1
X_26177_ _19935_/X _26177_/D vssd1 vssd1 vccd1 vccd1 _26177_/Q sky130_fd_sc_hd__dfxtp_1
X_23389_ _24759_/A _27243_/Q _27259_/Q _24804_/A _23388_/X vssd1 vssd1 vccd1 vccd1
+ _23393_/C sky130_fd_sc_hd__a221o_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13142_ _27287_/Q _13142_/B vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__and2_2
X_25128_ _27540_/Q _27519_/Q _18612_/B _25119_/X _18610_/X vssd1 vssd1 vccd1 vccd1
+ _25129_/B sky130_fd_sc_hd__a311o_1
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17950_ _27797_/Q _26558_/Q _26430_/Q _26110_/Q _17920_/X _17949_/X vssd1 vssd1 vccd1
+ vccd1 _17950_/X sky130_fd_sc_hd__mux4_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25059_ _27972_/A _25058_/X _25067_/S vssd1 vssd1 vccd1 vccd1 _25060_/A sky130_fd_sc_hd__mux2_1
X_13073_ _27062_/Q _13072_/X _13079_/S vssd1 vssd1 vccd1 vccd1 _13074_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16901_ _16897_/X _16898_/Y _16900_/Y vssd1 vssd1 vccd1 vccd1 _24264_/A sky130_fd_sc_hd__o21a_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17881_ _24624_/B _17881_/B _17881_/C vssd1 vssd1 vccd1 vccd1 _17882_/A sky130_fd_sc_hd__and3_1
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19620_ _19620_/A vssd1 vssd1 vccd1 vccd1 _19620_/X sky130_fd_sc_hd__clkbuf_1
X_16832_ _16800_/B _16830_/Y _16831_/Y vssd1 vssd1 vccd1 vccd1 _16832_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19551_ _26969_/Q _26937_/Q _26905_/Q _26873_/Q _19061_/X _18920_/X vssd1 vssd1 vccd1
+ vccd1 _19551_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16763_ _16752_/A _16754_/Y _16843_/A _16762_/Y vssd1 vssd1 vccd1 vccd1 _16763_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_13975_ _26802_/Q _13969_/X _13965_/X _13974_/Y vssd1 vssd1 vccd1 vccd1 _26802_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18502_ _18502_/A _18479_/X vssd1 vssd1 vccd1 vccd1 _18502_/X sky130_fd_sc_hd__or2b_1
X_15714_ _15714_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15714_/Y sky130_fd_sc_hd__nor2_1
XFILLER_202_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12926_ input44/X input45/X input46/X input47/X vssd1 vssd1 vccd1 vccd1 _12928_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19482_ _19482_/A vssd1 vssd1 vccd1 vccd1 _19482_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16694_ _16778_/A _16470_/A _16693_/X vssd1 vssd1 vccd1 vccd1 _16694_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18433_ _18379_/X _18430_/X _18432_/X _18384_/X vssd1 vssd1 vccd1 vccd1 _18433_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15645_ _13111_/X _26160_/Q _15645_/S vssd1 vssd1 vccd1 vccd1 _15646_/A sky130_fd_sc_hd__mux2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _18311_/X _18357_/X _18363_/X _18253_/X vssd1 vssd1 vccd1 vccd1 _18374_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_187_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15576_ _26191_/Q _14743_/A _15584_/S vssd1 vssd1 vccd1 vccd1 _15577_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17315_ _25937_/Q _26003_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17316_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14527_ _14527_/A vssd1 vssd1 vccd1 vccd1 _15779_/A sky130_fd_sc_hd__buf_2
X_18295_ _17912_/X _18294_/X _17915_/X vssd1 vssd1 vccd1 vccd1 _18295_/X sky130_fd_sc_hd__o21a_1
XFILLER_175_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17246_ _17307_/A vssd1 vssd1 vccd1 vccd1 _17295_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14458_ _26639_/Q _14441_/X _14455_/X _14457_/Y vssd1 vssd1 vccd1 vccd1 _26639_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_31_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _26974_/Q _13408_/X _13415_/S vssd1 vssd1 vccd1 vccd1 _13410_/A sky130_fd_sc_hd__mux2_1
X_14389_ _26660_/Q _14379_/X _14385_/X _14388_/Y vssd1 vssd1 vccd1 vccd1 _26660_/D
+ sky130_fd_sc_hd__a31o_1
X_17177_ _17299_/A vssd1 vssd1 vccd1 vccd1 _17177_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16128_ _16126_/Y _16119_/X _16121_/X _14425_/A _16127_/Y vssd1 vssd1 vccd1 vccd1
+ _24308_/A sky130_fd_sc_hd__o221a_1
XFILLER_115_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16059_ _27478_/Q _27270_/Q vssd1 vssd1 vccd1 vccd1 _16059_/X sky130_fd_sc_hd__and2_1
XFILLER_170_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19818_ _25726_/A vssd1 vssd1 vccd1 vccd1 _19887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19749_ _19814_/A vssd1 vssd1 vccd1 vccd1 _19749_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22760_ _22760_/A vssd1 vssd1 vccd1 vccd1 _22760_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21711_ _21705_/X _21706_/X _21707_/X _21708_/X _21709_/X _21710_/X vssd1 vssd1 vccd1
+ vccd1 _21712_/A sky130_fd_sc_hd__mux4_1
XFILLER_53_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22691_ _22681_/X _22682_/X _22683_/X _22684_/X _22685_/X _22686_/X vssd1 vssd1 vccd1
+ vccd1 _22692_/A sky130_fd_sc_hd__mux4_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24430_ _24430_/A vssd1 vssd1 vccd1 vccd1 _27493_/D sky130_fd_sc_hd__clkbuf_1
X_21642_ _21642_/A vssd1 vssd1 vccd1 vccd1 _21642_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24361_ _27563_/Q _24361_/B vssd1 vssd1 vccd1 vccd1 _24362_/A sky130_fd_sc_hd__and2_1
XANTENNA_20 _25996_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21573_ _21561_/X _21562_/X _21563_/X _21564_/X _21566_/X _21568_/X vssd1 vssd1 vccd1
+ vccd1 _21574_/A sky130_fd_sc_hd__mux4_1
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_31 _27838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26100_ _19669_/X _26100_/D vssd1 vssd1 vccd1 vccd1 _26100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23312_ _27742_/Q vssd1 vssd1 vccd1 vccd1 _23312_/Y sky130_fd_sc_hd__inv_2
XANTENNA_42 _18358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_53 _18134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27080_ _27112_/CLK _27080_/D vssd1 vssd1 vccd1 vccd1 _27080_/Q sky130_fd_sc_hd__dfxtp_1
X_20524_ _20512_/X _20513_/X _20514_/X _20515_/X _20517_/X _20519_/X vssd1 vssd1 vccd1
+ vccd1 _20525_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_64 _18312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24292_ _24304_/A vssd1 vssd1 vccd1 vccd1 _24302_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_75 _18493_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26031_ _27088_/CLK _26031_/D vssd1 vssd1 vccd1 vccd1 _26031_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_86 _24405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23243_ _23243_/A vssd1 vssd1 vccd1 vccd1 _27156_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_97 _19215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20455_ _20455_/A vssd1 vssd1 vccd1 vccd1 _20455_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23174_ _27126_/Q _17766_/X _23176_/S vssd1 vssd1 vccd1 vccd1 _23175_/A sky130_fd_sc_hd__mux2_1
X_20386_ _20376_/X _20377_/X _20378_/X _20379_/X _20380_/X _20381_/X vssd1 vssd1 vccd1
+ vccd1 _20387_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22125_ _22173_/A vssd1 vssd1 vccd1 vccd1 _22125_/X sky130_fd_sc_hd__clkbuf_1
X_27982_ _27982_/A _15902_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
XFILLER_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_713 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22056_ _22072_/A vssd1 vssd1 vccd1 vccd1 _22056_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26933_ _22574_/X _26933_/D vssd1 vssd1 vccd1 vccd1 _26933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21007_ _21039_/A vssd1 vssd1 vccd1 vccd1 _21007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26864_ _22330_/X _26864_/D vssd1 vssd1 vccd1 vccd1 _26864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25815_ _26014_/CLK _25815_/D vssd1 vssd1 vccd1 vccd1 _25815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26795_ _22092_/X _26795_/D vssd1 vssd1 vccd1 vccd1 _26795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13760_ _26874_/Q _13750_/X _13683_/B _13759_/Y vssd1 vssd1 vccd1 vccd1 _26874_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22958_ _22958_/A vssd1 vssd1 vccd1 vccd1 _22958_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25746_ _17437_/X _27830_/Q _25746_/S vssd1 vssd1 vccd1 vccd1 _25747_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21909_ _21895_/X _21896_/X _21897_/X _21898_/X _21899_/X _21900_/X vssd1 vssd1 vccd1
+ vccd1 _21910_/A sky130_fd_sc_hd__mux4_1
X_13691_ _13691_/A vssd1 vssd1 vccd1 vccd1 _13745_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25677_ _25709_/A vssd1 vssd1 vccd1 vccd1 _25677_/X sky130_fd_sc_hd__clkbuf_2
X_22889_ _22889_/A vssd1 vssd1 vccd1 vccd1 _22956_/A sky130_fd_sc_hd__buf_2
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15430_ _15430_/A vssd1 vssd1 vccd1 vccd1 _26256_/D sky130_fd_sc_hd__clkbuf_1
X_27416_ _27416_/CLK _27416_/D vssd1 vssd1 vccd1 vccd1 _27416_/Q sky130_fd_sc_hd__dfxtp_1
X_24628_ _16982_/C _24631_/B _24638_/B _24499_/X vssd1 vssd1 vccd1 vccd1 _27572_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_102_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15361_ _15361_/A vssd1 vssd1 vccd1 vccd1 _26287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24559_ _27641_/Q _24565_/B vssd1 vssd1 vccd1 vccd1 _24560_/A sky130_fd_sc_hd__and2_1
X_27347_ _27450_/CLK _27347_/D vssd1 vssd1 vccd1 vccd1 _27347_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17100_ _17052_/X _17093_/X _17096_/X _17099_/X vssd1 vssd1 vccd1 vccd1 _17100_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_184_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14312_ _14399_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14312_/Y sky130_fd_sc_hd__nor2_1
X_18080_ _26947_/Q _26915_/Q _26883_/Q _26851_/Q _17999_/X _18000_/X vssd1 vssd1 vccd1
+ vccd1 _18080_/X sky130_fd_sc_hd__mux4_2
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15292_ _15292_/A vssd1 vssd1 vccd1 vccd1 _26317_/D sky130_fd_sc_hd__clkbuf_1
X_27278_ _27278_/CLK _27278_/D vssd1 vssd1 vccd1 vccd1 _27278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14243_ _14257_/A vssd1 vssd1 vccd1 vccd1 _14248_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _17029_/X _17031_/B vssd1 vssd1 vccd1 vccd1 _17031_/X sky130_fd_sc_hd__and2b_1
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26229_ _20113_/X _26229_/D vssd1 vssd1 vccd1 vccd1 _26229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14174_ _14350_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14174_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ _27290_/Q _13125_/B vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__and2_1
XFILLER_98_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18982_ _19399_/A vssd1 vssd1 vccd1 vccd1 _18982_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _17779_/X _17926_/X _17931_/X _17932_/X vssd1 vssd1 vccd1 vccd1 _17947_/B
+ sky130_fd_sc_hd__a211o_1
X_13056_ _27301_/Q _13109_/B vssd1 vssd1 vccd1 vccd1 _13056_/X sky130_fd_sc_hd__and2_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater107 _27092_/CLK vssd1 vssd1 vccd1 vccd1 _25900_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_61_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17864_ _26811_/Q _26779_/Q _26747_/Q _26715_/Q _17863_/X _17805_/X vssd1 vssd1 vccd1
+ vccd1 _17864_/X sky130_fd_sc_hd__mux4_1
Xrepeater118 _27285_/CLK vssd1 vssd1 vccd1 vccd1 _27684_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater129 _26039_/CLK vssd1 vssd1 vccd1 vccd1 _26038_/CLK sky130_fd_sc_hd__clkbuf_1
X_19603_ _19589_/X _19590_/X _19591_/X _19592_/X _19593_/X _19594_/X vssd1 vssd1 vccd1
+ vccd1 _19604_/A sky130_fd_sc_hd__mux4_1
XFILLER_93_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _16815_/A _16815_/B vssd1 vssd1 vccd1 vccd1 _16815_/X sky130_fd_sc_hd__or2_1
XFILLER_4_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17795_ _18395_/A vssd1 vssd1 vccd1 vccd1 _17886_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1042 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19534_ _19534_/A _19534_/B vssd1 vssd1 vccd1 vccd1 _19534_/X sky130_fd_sc_hd__or2_1
XFILLER_35_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16746_ _16765_/B _16764_/B _16764_/A vssd1 vssd1 vccd1 vccd1 _16746_/X sky130_fd_sc_hd__or3b_1
X_13958_ _14032_/A vssd1 vssd1 vccd1 vccd1 _13974_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19465_ _19465_/A vssd1 vssd1 vccd1 vccd1 _19465_/X sky130_fd_sc_hd__buf_2
XFILLER_35_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16677_ _16737_/A _16737_/C _16737_/B vssd1 vssd1 vccd1 vccd1 _16738_/B sky130_fd_sc_hd__a21o_1
X_13889_ _13889_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13889_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18416_ _26289_/Q _26257_/Q _26225_/Q _26193_/Q _18301_/X _18324_/X vssd1 vssd1 vccd1
+ vccd1 _18416_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _13058_/X _26168_/Q _15634_/S vssd1 vssd1 vccd1 vccd1 _15629_/A sky130_fd_sc_hd__mux2_1
X_19396_ _19419_/A _19396_/B vssd1 vssd1 vccd1 vccd1 _19396_/X sky130_fd_sc_hd__or2_1
XFILLER_194_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18347_ _18020_/A _18346_/X _18014_/A vssd1 vssd1 vccd1 vccd1 _18347_/X sky130_fd_sc_hd__o21a_1
XFILLER_175_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15559_ _15559_/A vssd1 vssd1 vccd1 vccd1 _26199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18278_ _18278_/A _18207_/X vssd1 vssd1 vccd1 vccd1 _18278_/X sky130_fd_sc_hd__or2b_1
XFILLER_147_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput40 la1_data_in[9] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_4
X_17229_ _17216_/X _17229_/B vssd1 vssd1 vccd1 vccd1 _17229_/X sky130_fd_sc_hd__and2b_1
Xinput51 la1_oenb[19] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_4
XFILLER_190_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput62 la1_oenb[29] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_4
Xinput73 user_clock2 vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20240_ _20232_/X _20233_/X _20234_/X _20235_/X _20236_/X _20237_/X vssd1 vssd1 vccd1
+ vccd1 _20241_/A sky130_fd_sc_hd__mux4_1
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20171_ _20171_/A vssd1 vssd1 vccd1 vccd1 _20171_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1067 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23930_ _25930_/Q _25996_/Q _25829_/Q _26028_/Q _23899_/X _23929_/X vssd1 vssd1 vccd1
+ vccd1 _23930_/X sky130_fd_sc_hd__mux4_1
XFILLER_69_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23861_ _23861_/A vssd1 vssd1 vccd1 vccd1 _23861_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25600_ _27717_/Q _25568_/X _25569_/X vssd1 vssd1 vccd1 vccd1 _25600_/Y sky130_fd_sc_hd__a21oi_1
X_22812_ _22812_/A vssd1 vssd1 vccd1 vccd1 _22812_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26580_ _21348_/X _26580_/D vssd1 vssd1 vccd1 vccd1 _26580_/Q sky130_fd_sc_hd__dfxtp_1
X_23792_ _23740_/X _23790_/X _23791_/X _23768_/X vssd1 vssd1 vccd1 vccd1 _27274_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25531_ _25517_/X _25522_/X _25523_/X _24899_/B _25524_/X vssd1 vssd1 vccd1 vccd1
+ _25531_/X sky130_fd_sc_hd__o311a_1
X_22743_ _22735_/X _22736_/X _22737_/X _22738_/X _22739_/X _22740_/X vssd1 vssd1 vccd1
+ vccd1 _22744_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25462_ _25553_/A vssd1 vssd1 vccd1 vccd1 _25462_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22674_ _22674_/A vssd1 vssd1 vccd1 vccd1 _22674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_729 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24413_ _24538_/A vssd1 vssd1 vccd1 vccd1 _24422_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_27201_ _27352_/CLK _27201_/D vssd1 vssd1 vccd1 vccd1 _27201_/Q sky130_fd_sc_hd__dfxtp_1
X_21625_ _21615_/X _21616_/X _21617_/X _21618_/X _21619_/X _21620_/X vssd1 vssd1 vccd1
+ vccd1 _21626_/A sky130_fd_sc_hd__mux4_1
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25393_ _25415_/A vssd1 vssd1 vccd1 vccd1 _25402_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24344_ _27555_/Q _24350_/B vssd1 vssd1 vccd1 vccd1 _24345_/A sky130_fd_sc_hd__and2_1
X_27132_ _27132_/CLK _27132_/D vssd1 vssd1 vccd1 vccd1 _27132_/Q sky130_fd_sc_hd__dfxtp_1
X_21556_ _21556_/A vssd1 vssd1 vccd1 vccd1 _21556_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20507_ _20507_/A vssd1 vssd1 vccd1 vccd1 _20507_/X sky130_fd_sc_hd__clkbuf_1
X_27063_ _23022_/X _27063_/D vssd1 vssd1 vccd1 vccd1 _27063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24275_ _16215_/X _16217_/Y _16218_/X _24273_/X vssd1 vssd1 vccd1 vccd1 _27412_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21487_ _21475_/X _21476_/X _21477_/X _21478_/X _21480_/X _21482_/X vssd1 vssd1 vccd1
+ vccd1 _21488_/A sky130_fd_sc_hd__mux4_1
XFILLER_180_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26014_ _26014_/CLK _26014_/D vssd1 vssd1 vccd1 vccd1 _26014_/Q sky130_fd_sc_hd__dfxtp_1
X_23226_ _17485_/X _27149_/Q _23226_/S vssd1 vssd1 vccd1 vccd1 _23227_/A sky130_fd_sc_hd__mux2_1
X_20438_ _20424_/X _20425_/X _20426_/X _20427_/X _20430_/X _20433_/X vssd1 vssd1 vccd1
+ vccd1 _20439_/A sky130_fd_sc_hd__mux4_1
XFILLER_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23157_ _27118_/Q _17740_/X _23165_/S vssd1 vssd1 vccd1 vccd1 _23158_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20369_ _20369_/A vssd1 vssd1 vccd1 vccd1 _20369_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22108_ _22455_/A vssd1 vssd1 vccd1 vccd1 _22175_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23088_ _27088_/Q _17747_/X _23092_/S vssd1 vssd1 vccd1 vccd1 _23089_/A sky130_fd_sc_hd__mux2_1
X_27965_ _27965_/A _15911_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_88_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22039_ _22071_/A vssd1 vssd1 vccd1 vccd1 _22039_/X sky130_fd_sc_hd__clkbuf_2
X_26916_ _22512_/X _26916_/D vssd1 vssd1 vccd1 vccd1 _26916_/Q sky130_fd_sc_hd__dfxtp_1
X_14930_ _14930_/A vssd1 vssd1 vccd1 vccd1 _26470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26847_ _22274_/X _26847_/D vssd1 vssd1 vccd1 vccd1 _26847_/Q sky130_fd_sc_hd__dfxtp_1
X_14861_ _14861_/A vssd1 vssd1 vccd1 vccd1 _26501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16600_ _16879_/A _16879_/B _16878_/B _16902_/B _16599_/Y vssd1 vssd1 vccd1 vccd1
+ _16600_/Y sky130_fd_sc_hd__a311oi_2
X_13812_ _13904_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13812_/Y sky130_fd_sc_hd__nor2_1
X_17580_ _17495_/X _25865_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17581_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26778_ _22032_/X _26778_/D vssd1 vssd1 vccd1 vccd1 _26778_/Q sky130_fd_sc_hd__dfxtp_1
X_14792_ _14792_/A vssd1 vssd1 vccd1 vccd1 _14805_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16531_ _16623_/C vssd1 vssd1 vccd1 vccd1 _16535_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13743_ _13923_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13743_/Y sky130_fd_sc_hd__nor2_1
X_25729_ _25721_/X _25722_/X _25723_/X _25724_/X _25725_/X _25726_/X vssd1 vssd1 vccd1
+ vccd1 _25730_/A sky130_fd_sc_hd__mux4_1
XFILLER_188_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19250_ _19250_/A _19250_/B vssd1 vssd1 vccd1 vccd1 _19250_/X sky130_fd_sc_hd__or2_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16462_ _16778_/A _16462_/B vssd1 vssd1 vccd1 vccd1 _16471_/B sky130_fd_sc_hd__xnor2_1
XFILLER_189_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ _13762_/B _15190_/A vssd1 vssd1 vccd1 vccd1 _13691_/A sky130_fd_sc_hd__or2_1
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18201_ _26696_/Q _26664_/Q _26632_/Q _26600_/Q _18177_/X _18106_/X vssd1 vssd1 vccd1
+ vccd1 _18202_/A sky130_fd_sc_hd__mux4_1
XFILLER_19_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15413_ _15413_/A vssd1 vssd1 vccd1 vccd1 _26264_/D sky130_fd_sc_hd__clkbuf_1
X_19181_ _19158_/X _19180_/X _19089_/X vssd1 vssd1 vccd1 vccd1 _19181_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16393_ _16742_/A _16393_/B vssd1 vssd1 vccd1 vccd1 _16393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18132_ _26821_/Q _26789_/Q _26757_/Q _26725_/Q _18034_/X _18058_/X vssd1 vssd1 vccd1
+ vccd1 _18132_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15344_ _14721_/X _26294_/Q _15346_/S vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18063_ _18057_/X _18059_/X _18061_/X _18062_/X vssd1 vssd1 vccd1 vccd1 _18063_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15275_ _15332_/S vssd1 vssd1 vccd1 vccd1 _15284_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17014_ input35/X vssd1 vssd1 vccd1 vccd1 _17291_/A sky130_fd_sc_hd__buf_2
X_14226_ _14403_/A _14226_/B vssd1 vssd1 vccd1 vccd1 _14226_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ _14157_/A vssd1 vssd1 vccd1 vccd1 _14157_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13108_/A vssd1 vssd1 vccd1 vccd1 _13108_/X sky130_fd_sc_hd__buf_4
X_14088_ _14354_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14088_/Y sky130_fd_sc_hd__nor2_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ _18989_/A _18965_/B _18965_/C vssd1 vssd1 vccd1 vccd1 _18966_/A sky130_fd_sc_hd__and3_1
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _17912_/X _17914_/X _17915_/X vssd1 vssd1 vccd1 vccd1 _17916_/X sky130_fd_sc_hd__o21a_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _27269_/Q vssd1 vssd1 vccd1 vccd1 _16017_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18896_ _19401_/A vssd1 vssd1 vccd1 vccd1 _18896_/X sky130_fd_sc_hd__buf_4
XFILLER_79_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17847_ _17900_/A vssd1 vssd1 vccd1 vccd1 _18418_/A sky130_fd_sc_hd__buf_2
XFILLER_187_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17778_ _18443_/A vssd1 vssd1 vccd1 vccd1 _18150_/A sky130_fd_sc_hd__clkbuf_2
X_19517_ _26711_/Q _26679_/Q _26647_/Q _26615_/Q _18816_/X _18818_/X vssd1 vssd1 vccd1
+ vccd1 _19517_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16729_ _16076_/A _16767_/A _16450_/A _16084_/A vssd1 vssd1 vccd1 vccd1 _16729_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19448_ _19448_/A vssd1 vssd1 vccd1 vccd1 _19448_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19379_ _18814_/X _19378_/X _18785_/X vssd1 vssd1 vccd1 vccd1 _19379_/X sky130_fd_sc_hd__o21a_1
X_21410_ _21476_/A vssd1 vssd1 vccd1 vccd1 _21410_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22390_ _22422_/A vssd1 vssd1 vccd1 vccd1 _22390_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21341_ _21389_/A vssd1 vssd1 vccd1 vccd1 _21341_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24060_ _24060_/A vssd1 vssd1 vccd1 vccd1 _27307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21272_ _21304_/A vssd1 vssd1 vccd1 vccd1 _21272_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23011_ _25637_/A vssd1 vssd1 vccd1 vccd1 _23011_/X sky130_fd_sc_hd__clkbuf_1
X_20223_ _20223_/A vssd1 vssd1 vccd1 vccd1 _20223_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20154_ _20146_/X _20147_/X _20148_/X _20149_/X _20150_/X _20151_/X vssd1 vssd1 vccd1
+ vccd1 _20155_/A sky130_fd_sc_hd__mux4_1
XFILLER_44_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27750_ _27750_/CLK _27750_/D vssd1 vssd1 vccd1 vccd1 _27750_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20085_ _20085_/A vssd1 vssd1 vccd1 vccd1 _20085_/X sky130_fd_sc_hd__clkbuf_1
X_24962_ _24962_/A _24962_/B vssd1 vssd1 vccd1 vccd1 _24962_/Y sky130_fd_sc_hd__nand2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26701_ _21770_/X _26701_/D vssd1 vssd1 vccd1 vccd1 _26701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23913_ _27842_/Q _27146_/Q _25891_/Q _25859_/Q _23873_/X _23897_/X vssd1 vssd1 vccd1
+ vccd1 _23913_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27681_ _27681_/CLK _27681_/D vssd1 vssd1 vccd1 vccd1 _27972_/A sky130_fd_sc_hd__dfxtp_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24893_ _24893_/A _24896_/C vssd1 vssd1 vccd1 vccd1 _24894_/B sky130_fd_sc_hd__xnor2_1
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26632_ _21524_/X _26632_/D vssd1 vssd1 vccd1 vccd1 _26632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23844_ _23842_/X _23843_/X _23844_/S vssd1 vssd1 vccd1 vccd1 _23844_/X sky130_fd_sc_hd__mux2_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26563_ _21282_/X _26563_/D vssd1 vssd1 vccd1 vccd1 _26563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23775_ _27067_/Q _23761_/X _23763_/X _27099_/Q _23765_/X vssd1 vssd1 vccd1 vccd1
+ _23775_/X sky130_fd_sc_hd__a221o_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20987_ _20972_/X _20974_/X _20976_/X _20978_/X _20979_/X _20980_/X vssd1 vssd1 vccd1
+ vccd1 _20988_/A sky130_fd_sc_hd__mux4_1
XFILLER_41_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25514_ _25500_/X _25213_/B _25512_/X _25513_/X vssd1 vssd1 vccd1 vccd1 _25514_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22726_ _22726_/A vssd1 vssd1 vccd1 vccd1 _22726_/X sky130_fd_sc_hd__clkbuf_1
X_26494_ _21038_/X _26494_/D vssd1 vssd1 vccd1 vccd1 _26494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22657_ _22649_/X _22650_/X _22651_/X _22652_/X _22653_/X _22654_/X vssd1 vssd1 vccd1
+ vccd1 _22658_/A sky130_fd_sc_hd__mux4_1
XFILLER_139_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25445_ _27753_/Q _25437_/A _25110_/B _25625_/S vssd1 vssd1 vccd1 vccd1 _25466_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_186_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21608_ _21608_/A vssd1 vssd1 vccd1 vccd1 _21608_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13390_ _26980_/Q _13389_/X _13399_/S vssd1 vssd1 vccd1 vccd1 _13391_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22588_ _22588_/A vssd1 vssd1 vccd1 vccd1 _22588_/X sky130_fd_sc_hd__clkbuf_1
X_25376_ _27728_/Q input70/X _25380_/S vssd1 vssd1 vccd1 vccd1 _25377_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27115_ _27115_/CLK _27115_/D vssd1 vssd1 vccd1 vccd1 _27115_/Q sky130_fd_sc_hd__dfxtp_1
X_21539_ _21529_/X _21530_/X _21531_/X _21532_/X _21533_/X _21534_/X vssd1 vssd1 vccd1
+ vccd1 _21540_/A sky130_fd_sc_hd__mux4_1
XFILLER_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24327_ _24327_/A vssd1 vssd1 vccd1 vccd1 _27447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_794 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15060_ _14727_/X _26420_/Q _15068_/S vssd1 vssd1 vccd1 vccd1 _15061_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24258_ _24258_/A _24264_/B vssd1 vssd1 vccd1 vccd1 _27401_/D sky130_fd_sc_hd__nor2_1
X_27046_ _22966_/X _27046_/D vssd1 vssd1 vccd1 vccd1 _27046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14011_ _26792_/Q _14005_/X _14001_/X _14010_/Y vssd1 vssd1 vccd1 vccd1 _26792_/D
+ sky130_fd_sc_hd__a31o_1
X_23209_ _17460_/X _27141_/Q _23215_/S vssd1 vssd1 vccd1 vccd1 _23210_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24189_ _27470_/Q _24195_/B vssd1 vssd1 vccd1 vccd1 _24190_/A sky130_fd_sc_hd__and2_1
XFILLER_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_874 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18750_ _18750_/A vssd1 vssd1 vccd1 vccd1 _26035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15962_ _15980_/A vssd1 vssd1 vccd1 vccd1 _15967_/A sky130_fd_sc_hd__buf_2
X_27948_ _27948_/A _15987_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17701_ _17701_/A vssd1 vssd1 vccd1 vccd1 _25919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14913_ _14913_/A vssd1 vssd1 vccd1 vccd1 _26478_/D sky130_fd_sc_hd__clkbuf_1
X_18681_ _26005_/Q _17763_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _18682_/A sky130_fd_sc_hd__mux2_1
X_15893_ _15893_/A vssd1 vssd1 vccd1 vccd1 _15893_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17632_ _17466_/X _25888_/Q _17634_/S vssd1 vssd1 vccd1 vccd1 _17633_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14844_ _26508_/Q _13363_/X _14846_/S vssd1 vssd1 vccd1 vccd1 _14845_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17563_ _17563_/A vssd1 vssd1 vccd1 vccd1 _25857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14775_ _14775_/A vssd1 vssd1 vccd1 vccd1 _14775_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19302_ _18895_/A _19296_/X _19299_/X _19301_/X vssd1 vssd1 vccd1 vccd1 _19302_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _16672_/A _16700_/B _16631_/A _16664_/A vssd1 vssd1 vccd1 vccd1 _16514_/X
+ sky130_fd_sc_hd__and4_1
X_13726_ _26888_/Q _13724_/X _13718_/X _13725_/Y vssd1 vssd1 vccd1 vccd1 _26888_/D
+ sky130_fd_sc_hd__a31o_1
X_17494_ _17494_/A vssd1 vssd1 vccd1 vccd1 _25832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19233_ _19391_/A vssd1 vssd1 vccd1 vccd1 _19346_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ _16445_/A _16445_/B vssd1 vssd1 vccd1 vccd1 _16445_/X sky130_fd_sc_hd__or2_1
X_13657_ _13926_/A _13661_/B vssd1 vssd1 vccd1 vccd1 _13657_/Y sky130_fd_sc_hd__nor2_1
X_19164_ _19157_/X _19160_/X _19163_/X _19022_/X _19139_/X vssd1 vssd1 vccd1 vccd1
+ _19175_/B sky130_fd_sc_hd__a221o_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _23035_/A _16508_/B _16536_/B _14507_/A _16375_/Y vssd1 vssd1 vccd1 vccd1
+ _16749_/B sky130_fd_sc_hd__o221a_1
XFILLER_185_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13588_ _13602_/A vssd1 vssd1 vccd1 vccd1 _13593_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18115_ _26276_/Q _26244_/Q _26212_/Q _26180_/Q _18044_/X _18068_/X vssd1 vssd1 vccd1
+ vccd1 _18115_/X sky130_fd_sc_hd__mux4_2
XFILLER_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15327_ _15327_/A vssd1 vssd1 vccd1 vccd1 _26301_/D sky130_fd_sc_hd__clkbuf_1
X_19095_ _19086_/X _19090_/X _19094_/X _19022_/X _19023_/X vssd1 vssd1 vccd1 vccd1
+ _19107_/B sky130_fd_sc_hd__a221o_1
XFILLER_9_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18046_ _18020_/X _18045_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _18046_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ _14807_/X _26331_/Q _15260_/S vssd1 vssd1 vccd1 vccd1 _15259_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14209_ _26725_/Q _14199_/X _14207_/X _14208_/Y vssd1 vssd1 vccd1 vccd1 _26725_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _15189_/A vssd1 vssd1 vccd1 vccd1 _26362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19997_ _20065_/A vssd1 vssd1 vccd1 vccd1 _19997_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18948_ _18938_/X _18942_/X _18947_/X _18854_/X _18880_/X vssd1 vssd1 vccd1 vccd1
+ _18965_/B sky130_fd_sc_hd__a221o_1
XFILLER_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18879_ _27602_/Q vssd1 vssd1 vccd1 vccd1 _19393_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20910_ _20942_/A vssd1 vssd1 vccd1 vccd1 _20910_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21890_ _21890_/A vssd1 vssd1 vccd1 vccd1 _21890_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20841_ _20841_/A vssd1 vssd1 vccd1 vccd1 _20841_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23560_ _23560_/A _23560_/B vssd1 vssd1 vccd1 vccd1 _23561_/A sky130_fd_sc_hd__and2_1
X_20772_ _20772_/A vssd1 vssd1 vccd1 vccd1 _20772_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22511_ _22503_/X _22504_/X _22505_/X _22506_/X _22507_/X _22508_/X vssd1 vssd1 vccd1
+ vccd1 _22512_/A sky130_fd_sc_hd__mux4_1
XFILLER_50_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23491_ _27189_/Q _23495_/B vssd1 vssd1 vccd1 vccd1 _23491_/X sky130_fd_sc_hd__or2_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22442_ _22442_/A vssd1 vssd1 vccd1 vccd1 _22442_/X sky130_fd_sc_hd__clkbuf_1
X_25230_ _25261_/A _25230_/B vssd1 vssd1 vccd1 vccd1 _25230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25161_ _27526_/Q _27494_/Q vssd1 vssd1 vccd1 vccd1 _25162_/B sky130_fd_sc_hd__or2_1
X_22373_ _22421_/A vssd1 vssd1 vccd1 vccd1 _22373_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24112_ _24112_/A vssd1 vssd1 vccd1 vccd1 _27330_/D sky130_fd_sc_hd__clkbuf_1
X_21324_ _21390_/A vssd1 vssd1 vccd1 vccd1 _21324_/X sky130_fd_sc_hd__clkbuf_1
X_25092_ _27840_/Q _27144_/Q _25889_/Q _25857_/Q _25061_/X _24975_/X vssd1 vssd1 vccd1
+ vccd1 _25092_/X sky130_fd_sc_hd__mux4_1
XFILLER_191_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24043_ _27857_/Q _27161_/Q _25906_/Q _25874_/Q _24014_/X _23749_/X vssd1 vssd1 vccd1
+ vccd1 _24043_/X sky130_fd_sc_hd__mux4_1
X_21255_ _21303_/A vssd1 vssd1 vccd1 vccd1 _21255_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20206_ _20200_/X _20201_/X _20202_/X _20203_/X _20204_/X _20205_/X vssd1 vssd1 vccd1
+ vccd1 _20207_/A sky130_fd_sc_hd__mux4_1
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21186_ _21186_/A vssd1 vssd1 vccd1 vccd1 _21186_/X sky130_fd_sc_hd__clkbuf_1
X_27802_ _25664_/X _27802_/D vssd1 vssd1 vccd1 vccd1 _27802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20137_ _20137_/A vssd1 vssd1 vccd1 vccd1 _20137_/X sky130_fd_sc_hd__clkbuf_1
X_25994_ _25995_/CLK _25994_/D vssd1 vssd1 vccd1 vccd1 _25994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27733_ _27737_/CLK _27733_/D vssd1 vssd1 vccd1 vccd1 _27733_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ _20060_/X _20061_/X _20062_/X _20063_/X _20064_/X _20065_/X vssd1 vssd1 vccd1
+ vccd1 _20069_/A sky130_fd_sc_hd__mux4_1
XFILLER_57_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24945_ _27665_/Q _24935_/X _24944_/Y _24938_/X vssd1 vssd1 vccd1 vccd1 _27665_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27664_ _27666_/CLK _27664_/D vssd1 vssd1 vccd1 vccd1 _27664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24876_ _27651_/Q _24861_/X _24875_/Y _24864_/X vssd1 vssd1 vccd1 vccd1 _27651_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 _27356_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater290 _27357_/CLK vssd1 vssd1 vccd1 vccd1 _27335_/CLK sky130_fd_sc_hd__clkbuf_1
X_26615_ _21466_/X _26615_/D vssd1 vssd1 vccd1 vccd1 _26615_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 _18396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 _19276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23827_ _27833_/Q _27137_/Q _25882_/Q _25850_/Q _23826_/X _23802_/X vssd1 vssd1 vccd1
+ vccd1 _23827_/X sky130_fd_sc_hd__mux4_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27595_ _27601_/CLK _27595_/D vssd1 vssd1 vccd1 vccd1 _27595_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 _13166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _13417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_357 _14724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14560_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14571_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_368 _27859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26546_ _21222_/X _26546_/D vssd1 vssd1 vccd1 vccd1 _26546_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 _17950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23758_ _24047_/S vssd1 vssd1 vccd1 vccd1 _23797_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _27350_/Q _13108_/X _13102_/X _27318_/Q _13148_/X vssd1 vssd1 vccd1 vccd1
+ _16451_/A sky130_fd_sc_hd__a221oi_4
XFILLER_199_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22709_ _22697_/X _22698_/X _22699_/X _22700_/X _22702_/X _22704_/X vssd1 vssd1 vccd1
+ vccd1 _22710_/A sky130_fd_sc_hd__mux4_1
X_14491_ _26630_/Q _14478_/X _14474_/X _14490_/Y vssd1 vssd1 vccd1 vccd1 _26630_/D
+ sky130_fd_sc_hd__a31o_1
X_26477_ _20986_/X _26477_/D vssd1 vssd1 vccd1 vccd1 _26477_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23689_ _23689_/A vssd1 vssd1 vccd1 vccd1 _27249_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16230_/A _16235_/B _16240_/C vssd1 vssd1 vccd1 vccd1 _16230_/X sky130_fd_sc_hd__and3_1
X_13442_ _13861_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13442_/Y sky130_fd_sc_hd__nor2_1
X_25428_ _27752_/Q input65/X _25428_/S vssd1 vssd1 vccd1 vccd1 _25429_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13373_ _16252_/A vssd1 vssd1 vccd1 vccd1 _13373_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ _16249_/B vssd1 vssd1 vccd1 vccd1 _16276_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25359_ _25415_/A vssd1 vssd1 vccd1 vccd1 _25428_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ _14804_/X _26396_/Q _15112_/S vssd1 vssd1 vccd1 vccd1 _15113_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16092_ _16738_/A vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15043_ _15781_/A _15043_/B vssd1 vssd1 vccd1 vccd1 _15043_/Y sky130_fd_sc_hd__nor2_1
X_19920_ _20268_/A vssd1 vssd1 vccd1 vccd1 _19989_/A sky130_fd_sc_hd__clkbuf_2
X_27029_ _22906_/X _27029_/D vssd1 vssd1 vccd1 vccd1 _27029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19851_ _19899_/A vssd1 vssd1 vccd1 vccd1 _19851_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18802_ _27602_/Q vssd1 vssd1 vccd1 vccd1 _24407_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19782_ _19814_/A vssd1 vssd1 vccd1 vccd1 _19782_/X sky130_fd_sc_hd__clkbuf_1
X_16994_ _17325_/A vssd1 vssd1 vccd1 vccd1 _17382_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18733_ _26028_/Q _17734_/X _18735_/S vssd1 vssd1 vccd1 vccd1 _18734_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15945_ _15949_/A vssd1 vssd1 vccd1 vccd1 _15945_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18664_ _18664_/A vssd1 vssd1 vccd1 vccd1 _25997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _15894_/A vssd1 vssd1 vccd1 vccd1 _15881_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ _17440_/X _25880_/Q _17623_/S vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14827_ _26516_/Q _13337_/X _14835_/S vssd1 vssd1 vccd1 vccd1 _14828_/A sky130_fd_sc_hd__mux2_1
X_18595_ _27688_/Q vssd1 vssd1 vccd1 vccd1 _25568_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17546_ _17546_/A vssd1 vssd1 vccd1 vccd1 _25849_/D sky130_fd_sc_hd__clkbuf_1
X_14758_ _14758_/A vssd1 vssd1 vccd1 vccd1 _26539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ _26894_/Q _13697_/X _13705_/X _13708_/Y vssd1 vssd1 vccd1 vccd1 _26894_/D
+ sky130_fd_sc_hd__a31o_1
X_17477_ _17476_/X _25827_/Q _17486_/S vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14689_ _15762_/A _14699_/B vssd1 vssd1 vccd1 vccd1 _14689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19216_ _26153_/Q _26089_/Q _27017_/Q _26985_/Q _18807_/X _18810_/X vssd1 vssd1 vccd1
+ vccd1 _19217_/B sky130_fd_sc_hd__mux4_1
X_16428_ _16428_/A vssd1 vssd1 vccd1 vccd1 _16722_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19147_ _26406_/Q _26374_/Q _26342_/Q _26310_/Q _19054_/X _19100_/X vssd1 vssd1 vccd1
+ vccd1 _19147_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _16359_/A vssd1 vssd1 vccd1 vccd1 _16447_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_173_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19078_ _26403_/Q _26371_/Q _26339_/Q _26307_/Q _19054_/X _18982_/X vssd1 vssd1 vccd1
+ vccd1 _19078_/X sky130_fd_sc_hd__mux4_1
XFILLER_161_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18029_ _18029_/A vssd1 vssd1 vccd1 vccd1 _25950_/D sky130_fd_sc_hd__clkbuf_1
X_21040_ _21040_/A vssd1 vssd1 vccd1 vccd1 _21040_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22991_ _22974_/X _22976_/X _22978_/X _22980_/X _22981_/X _22982_/X vssd1 vssd1 vccd1
+ vccd1 _22992_/A sky130_fd_sc_hd__mux4_1
XFILLER_55_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24730_ _27608_/Q _24727_/X _24728_/X _24729_/X vssd1 vssd1 vccd1 vccd1 _27608_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21942_ _21942_/A vssd1 vssd1 vccd1 vccd1 _21942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21873_ _21863_/X _21864_/X _21865_/X _21866_/X _21867_/X _21868_/X vssd1 vssd1 vccd1
+ vccd1 _21874_/A sky130_fd_sc_hd__mux4_1
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24661_ _25540_/A vssd1 vssd1 vccd1 vccd1 _24671_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26400_ _20713_/X _26400_/D vssd1 vssd1 vccd1 vccd1 _26400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20824_ _20816_/X _20817_/X _20818_/X _20819_/X _20820_/X _20821_/X vssd1 vssd1 vccd1
+ vccd1 _20825_/A sky130_fd_sc_hd__mux4_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23612_ _25601_/A _27223_/Q _23616_/S vssd1 vssd1 vccd1 vccd1 _23613_/B sky130_fd_sc_hd__mux2_1
X_27380_ _27397_/CLK _27380_/D vssd1 vssd1 vccd1 vccd1 _27380_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24592_ _27656_/Q _24598_/B vssd1 vssd1 vccd1 vccd1 _24593_/A sky130_fd_sc_hd__and2_1
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26331_ _20473_/X _26331_/D vssd1 vssd1 vccd1 vccd1 _26331_/Q sky130_fd_sc_hd__dfxtp_1
X_20755_ _20771_/A vssd1 vssd1 vccd1 vccd1 _20755_/X sky130_fd_sc_hd__clkbuf_1
X_23543_ _23543_/A _23543_/B vssd1 vssd1 vccd1 vccd1 _23544_/A sky130_fd_sc_hd__and2_1
XFILLER_145_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23474_ _25132_/A vssd1 vssd1 vccd1 vccd1 _23474_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26262_ _20227_/X _26262_/D vssd1 vssd1 vccd1 vccd1 _26262_/Q sky130_fd_sc_hd__dfxtp_1
X_20686_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20686_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_28001_ _28001_/A _15879_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_195_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22425_ _22417_/X _22418_/X _22419_/X _22420_/X _22421_/X _22422_/X vssd1 vssd1 vccd1
+ vccd1 _22426_/A sky130_fd_sc_hd__mux4_1
X_25213_ _25221_/A _25213_/B vssd1 vssd1 vccd1 vccd1 _25213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26193_ _19985_/X _26193_/D vssd1 vssd1 vccd1 vccd1 _26193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22356_ _22356_/A vssd1 vssd1 vccd1 vccd1 _22356_/X sky130_fd_sc_hd__clkbuf_1
X_25144_ _25309_/A vssd1 vssd1 vccd1 vccd1 _25182_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21307_ _21377_/A vssd1 vssd1 vccd1 vccd1 _21307_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25075_ _25075_/A vssd1 vssd1 vccd1 vccd1 _25104_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22287_ _22335_/A vssd1 vssd1 vccd1 vccd1 _22287_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24026_ _24024_/X _24025_/X _24033_/S vssd1 vssd1 vccd1 vccd1 _24026_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21238_ _22546_/A vssd1 vssd1 vccd1 vccd1 _21585_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21169_ _21163_/X _21164_/X _21165_/X _21166_/X _21167_/X _21168_/X vssd1 vssd1 vccd1
+ vccd1 _21170_/A sky130_fd_sc_hd__mux4_1
XFILLER_46_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13991_ _14464_/A vssd1 vssd1 vccd1 vccd1 _14363_/A sky130_fd_sc_hd__buf_2
XFILLER_19_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25977_ _27783_/CLK _25977_/D vssd1 vssd1 vccd1 vccd1 _25977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15730_ _15730_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15730_/Y sky130_fd_sc_hd__nor2_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27716_ _27716_/CLK _27716_/D vssd1 vssd1 vccd1 vccd1 _27716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12942_ _23650_/A vssd1 vssd1 vccd1 vccd1 _23598_/A sky130_fd_sc_hd__buf_6
X_24928_ _24937_/A _24928_/B vssd1 vssd1 vccd1 vccd1 _24928_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27647_ _27667_/CLK _27647_/D vssd1 vssd1 vccd1 vccd1 _27647_/Q sky130_fd_sc_hd__dfxtp_1
X_15661_ _13150_/X _26153_/Q _15667_/S vssd1 vssd1 vccd1 vccd1 _15662_/A sky130_fd_sc_hd__mux2_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24859_ _24863_/A _24859_/B vssd1 vssd1 vccd1 vccd1 _24859_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_110 _19977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _22546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _25733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _25659_/A vssd1 vssd1 vccd1 vccd1 _19836_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14612_ _15775_/A _14620_/B vssd1 vssd1 vccd1 vccd1 _14612_/Y sky130_fd_sc_hd__nor2_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _13038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18380_ _18380_/A vssd1 vssd1 vccd1 vccd1 _18380_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15592_ _15592_/A vssd1 vssd1 vccd1 vccd1 _26184_/D sky130_fd_sc_hd__clkbuf_1
X_27578_ _27578_/CLK _27578_/D vssd1 vssd1 vccd1 vccd1 _27578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _13319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_165 _13398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _14452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17303_/X _17330_/X _17281_/X vssd1 vssd1 vccd1 vccd1 _17331_/X sky130_fd_sc_hd__a21bo_1
XANTENNA_187 _16495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _14493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14543_ _26615_/Q _14530_/X _14536_/X _14542_/Y vssd1 vssd1 vccd1 vccd1 _26615_/D
+ sky130_fd_sc_hd__a31o_1
X_26529_ _21162_/X _26529_/D vssd1 vssd1 vccd1 vccd1 _26529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17262_ _27215_/Q _17260_/X _17311_/S vssd1 vssd1 vccd1 vccd1 _17263_/A sky130_fd_sc_hd__mux2_1
X_14474_ _14510_/A vssd1 vssd1 vccd1 vccd1 _14474_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19001_ _18999_/X _19000_/X _19047_/S vssd1 vssd1 vccd1 vccd1 _19001_/X sky130_fd_sc_hd__mux2_1
X_16213_ _27525_/Q _15991_/A vssd1 vssd1 vccd1 vccd1 _16213_/X sky130_fd_sc_hd__or2b_1
XFILLER_186_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ _13425_/A _13672_/A _13672_/B vssd1 vssd1 vccd1 vccd1 _15623_/B sky130_fd_sc_hd__or3_2
XFILLER_186_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17193_ _25927_/Q _25993_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17194_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16144_ _27400_/Q _16144_/B vssd1 vssd1 vccd1 vccd1 _16144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13356_ _13356_/A vssd1 vssd1 vccd1 vccd1 _26991_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16075_ _16625_/A vssd1 vssd1 vccd1 vccd1 _16076_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13287_ _27016_/Q _13156_/X _13291_/S vssd1 vssd1 vccd1 vccd1 _13288_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ _15764_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15026_/Y sky130_fd_sc_hd__nor2_1
X_19903_ _19976_/A vssd1 vssd1 vccd1 vccd1 _19903_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19834_ _19834_/A vssd1 vssd1 vccd1 vccd1 _19900_/A sky130_fd_sc_hd__buf_2
XFILLER_151_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19765_ _19813_/A vssd1 vssd1 vccd1 vccd1 _19765_/X sky130_fd_sc_hd__clkbuf_1
X_16977_ _16977_/A vssd1 vssd1 vccd1 vccd1 _25910_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18716_ _26020_/Q _17708_/X _18724_/S vssd1 vssd1 vccd1 vccd1 _18717_/A sky130_fd_sc_hd__mux2_1
X_15928_ _15930_/A vssd1 vssd1 vccd1 vccd1 _15928_/Y sky130_fd_sc_hd__inv_2
X_19696_ _19728_/A vssd1 vssd1 vccd1 vccd1 _19696_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18647_ _18647_/A vssd1 vssd1 vccd1 vccd1 _25989_/D sky130_fd_sc_hd__clkbuf_1
X_15859_ _15862_/A vssd1 vssd1 vccd1 vccd1 _15859_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18578_ _26553_/Q _26521_/Q _26489_/Q _27065_/Q _17846_/X _17848_/X vssd1 vssd1 vccd1
+ vccd1 _18578_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17529_ _25735_/C _18691_/B vssd1 vssd1 vccd1 vccd1 _17586_/A sky130_fd_sc_hd__or2_4
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20540_ _20531_/X _20533_/X _20535_/X _20537_/X _20538_/X _20539_/X vssd1 vssd1 vccd1
+ vccd1 _20541_/A sky130_fd_sc_hd__mux4_1
X_20471_ _20471_/A vssd1 vssd1 vccd1 vccd1 _20471_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22210_ _22210_/A vssd1 vssd1 vccd1 vccd1 _22210_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23190_ _23190_/A vssd1 vssd1 vccd1 vccd1 _27132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22141_ _22173_/A vssd1 vssd1 vccd1 vccd1 _22141_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22072_ _22072_/A vssd1 vssd1 vccd1 vccd1 _22072_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25900_ _25900_/CLK _25900_/D vssd1 vssd1 vccd1 vccd1 _25900_/Q sky130_fd_sc_hd__dfxtp_1
X_21023_ _21039_/A vssd1 vssd1 vccd1 vccd1 _21023_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26880_ _22392_/X _26880_/D vssd1 vssd1 vccd1 vccd1 _26880_/Q sky130_fd_sc_hd__dfxtp_1
X_25831_ _26002_/CLK _25831_/D vssd1 vssd1 vccd1 vccd1 _25831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25762_ _17460_/X _27837_/Q _25768_/S vssd1 vssd1 vccd1 vccd1 _25763_/A sky130_fd_sc_hd__mux2_1
X_22974_ _25635_/A vssd1 vssd1 vccd1 vccd1 _22974_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27501_ _27623_/CLK _27501_/D vssd1 vssd1 vccd1 vccd1 _27501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24713_ _24841_/A vssd1 vssd1 vccd1 vccd1 _24771_/A sky130_fd_sc_hd__clkbuf_2
X_21925_ _21911_/X _21912_/X _21913_/X _21914_/X _21916_/X _21918_/X vssd1 vssd1 vccd1
+ vccd1 _21926_/A sky130_fd_sc_hd__mux4_1
X_25693_ _25709_/A vssd1 vssd1 vccd1 vccd1 _25693_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27432_ _27436_/CLK _27432_/D vssd1 vssd1 vccd1 vccd1 _27432_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24644_ _25434_/A vssd1 vssd1 vccd1 vccd1 _25540_/A sky130_fd_sc_hd__buf_2
X_21856_ _21856_/A vssd1 vssd1 vccd1 vccd1 _21856_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27363_ _27825_/CLK _27363_/D vssd1 vssd1 vccd1 vccd1 _27363_/Q sky130_fd_sc_hd__dfxtp_2
X_20807_ _20807_/A vssd1 vssd1 vccd1 vccd1 _20807_/X sky130_fd_sc_hd__clkbuf_1
X_21787_ _21777_/X _21778_/X _21779_/X _21780_/X _21781_/X _21782_/X vssd1 vssd1 vccd1
+ vccd1 _21788_/A sky130_fd_sc_hd__mux4_1
X_24575_ _24575_/A vssd1 vssd1 vccd1 vccd1 _27548_/D sky130_fd_sc_hd__clkbuf_1
X_26314_ _20407_/X _26314_/D vssd1 vssd1 vccd1 vccd1 _26314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23526_ _23526_/A _23526_/B vssd1 vssd1 vccd1 vccd1 _23527_/A sky130_fd_sc_hd__and2_1
XFILLER_168_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27294_ _27294_/CLK _27294_/D vssd1 vssd1 vccd1 vccd1 _27294_/Q sky130_fd_sc_hd__dfxtp_1
X_20738_ _20770_/A vssd1 vssd1 vccd1 vccd1 _20738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26245_ _20171_/X _26245_/D vssd1 vssd1 vccd1 vccd1 _26245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23457_ input14/X _23455_/X _23456_/X _23447_/X vssd1 vssd1 vccd1 vccd1 _27176_/D
+ sky130_fd_sc_hd__o211a_1
X_20669_ _20685_/A vssd1 vssd1 vccd1 vccd1 _20669_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13210_ _16224_/A vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22408_ _22408_/A vssd1 vssd1 vccd1 vccd1 _22408_/X sky130_fd_sc_hd__clkbuf_1
X_14190_ _14367_/A _14200_/B vssd1 vssd1 vccd1 vccd1 _14190_/Y sky130_fd_sc_hd__nor2_1
X_26176_ _19933_/X _26176_/D vssd1 vssd1 vccd1 vccd1 _26176_/Q sky130_fd_sc_hd__dfxtp_1
X_23388_ _24794_/A _27256_/Q _23333_/Y _27782_/Q vssd1 vssd1 vccd1 vccd1 _23388_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25127_ _25127_/A _25126_/X vssd1 vssd1 vccd1 vccd1 _25130_/A sky130_fd_sc_hd__or2b_1
X_13141_ _13141_/A vssd1 vssd1 vccd1 vccd1 _27051_/D sky130_fd_sc_hd__clkbuf_1
X_22339_ _22331_/X _22332_/X _22333_/X _22334_/X _22335_/X _22336_/X vssd1 vssd1 vccd1
+ vccd1 _22340_/A sky130_fd_sc_hd__mux4_1
XFILLER_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _14721_/A vssd1 vssd1 vccd1 vccd1 _13072_/X sky130_fd_sc_hd__buf_2
XFILLER_183_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25058_ _25055_/X _25057_/X _25074_/S vssd1 vssd1 vccd1 vccd1 _25058_/X sky130_fd_sc_hd__mux2_2
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16900_ _16308_/A _16790_/B _16899_/X vssd1 vssd1 vccd1 vccd1 _16900_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24009_ _24007_/X _24008_/X _24031_/S vssd1 vssd1 vccd1 vccd1 _24009_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17880_ _17872_/X _17875_/X _17879_/X _17854_/X _17856_/X vssd1 vssd1 vccd1 vccd1
+ _17881_/C sky130_fd_sc_hd__a221o_1
X_16831_ _16831_/A _16831_/B vssd1 vssd1 vccd1 vccd1 _16831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19550_ _19550_/A vssd1 vssd1 vccd1 vccd1 _26072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16762_ _16758_/Y _16842_/B _16761_/X vssd1 vssd1 vccd1 vccd1 _16762_/Y sky130_fd_sc_hd__a21oi_1
X_13974_ _14350_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _13974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_1174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18501_ _26165_/Q _26101_/Q _27029_/Q _26997_/Q _18455_/X _18011_/X vssd1 vssd1 vccd1
+ vccd1 _18502_/A sky130_fd_sc_hd__mux4_2
X_15713_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15713_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19481_ _19475_/X _19477_/X _19480_/X _18837_/X _19393_/X vssd1 vssd1 vccd1 vccd1
+ _19495_/B sky130_fd_sc_hd__a221o_1
XFILLER_111_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ input67/X input68/X input69/X input70/X vssd1 vssd1 vccd1 vccd1 _12928_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_74_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16693_ _16076_/A _16778_/A _16470_/A _16699_/A vssd1 vssd1 vccd1 vccd1 _16693_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18432_ _18432_/A _18317_/X vssd1 vssd1 vccd1 vccd1 _18432_/X sky130_fd_sc_hd__or2b_1
X_15644_ _15644_/A vssd1 vssd1 vccd1 vccd1 _26161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18198_/X _18359_/X _18362_/X _18203_/X vssd1 vssd1 vccd1 vccd1 _18363_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15621_/S vssd1 vssd1 vccd1 vccd1 _15584_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _27851_/Q _27155_/Q _25900_/Q _25868_/Q _17264_/X _17313_/X vssd1 vssd1 vccd1
+ vccd1 _17314_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _26620_/Q _14514_/X _14510_/X _14525_/Y vssd1 vssd1 vccd1 vccd1 _26620_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18294_ _26828_/Q _26796_/Q _26764_/Q _26732_/Q _18085_/X _17913_/X vssd1 vssd1 vccd1
+ vccd1 _18294_/X sky130_fd_sc_hd__mux4_2
X_17245_ _17238_/X _17239_/X _17241_/X _17244_/X vssd1 vssd1 vccd1 vccd1 _17245_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14457_ _15728_/A _14465_/B vssd1 vssd1 vccd1 vccd1 _14457_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13408_ _14798_/A vssd1 vssd1 vccd1 vccd1 _13408_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17176_ _17176_/A vssd1 vssd1 vccd1 vccd1 _27929_/A sky130_fd_sc_hd__clkbuf_1
X_14388_ _14388_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _14388_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16127_ _27405_/Q _16287_/A vssd1 vssd1 vccd1 vccd1 _16127_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13339_ _26996_/Q _13337_/X _13351_/S vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ _16052_/Y _16017_/B _16014_/B _16053_/Y vssd1 vssd1 vccd1 vccd1 _16063_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15009_ _26440_/Q _15002_/X _15003_/X _15008_/Y vssd1 vssd1 vccd1 vccd1 _26440_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19817_ _19886_/A vssd1 vssd1 vccd1 vccd1 _19817_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19748_ _19834_/A vssd1 vssd1 vccd1 vccd1 _19814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19679_ _19727_/A vssd1 vssd1 vccd1 vccd1 _19679_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21710_ _21726_/A vssd1 vssd1 vccd1 vccd1 _21710_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22690_ _22690_/A vssd1 vssd1 vccd1 vccd1 _22690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ _21631_/X _21632_/X _21633_/X _21634_/X _21635_/X _21636_/X vssd1 vssd1 vccd1
+ vccd1 _21642_/A sky130_fd_sc_hd__mux4_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21572_ _21572_/A vssd1 vssd1 vccd1 vccd1 _21572_/X sky130_fd_sc_hd__clkbuf_1
X_24360_ _24360_/A vssd1 vssd1 vccd1 vccd1 _27462_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_10 _25855_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _26024_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_32 _27840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23311_ _27726_/Q _23288_/Y _23262_/Y input59/X _23310_/Y vssd1 vssd1 vccd1 vccd1
+ _23320_/A sky130_fd_sc_hd__a221o_1
X_20523_ _20523_/A vssd1 vssd1 vccd1 vccd1 _20523_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_43 _17903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 _18202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24291_ _24291_/A vssd1 vssd1 vccd1 vccd1 _27423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_65 _18323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 _18516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26030_ _26030_/CLK _26030_/D vssd1 vssd1 vccd1 vccd1 _26030_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_87 _24405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23242_ _17508_/X _27156_/Q _23248_/S vssd1 vssd1 vccd1 vccd1 _23243_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_98 _19246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20454_ _20445_/X _20447_/X _20449_/X _20451_/X _20452_/X _20453_/X vssd1 vssd1 vccd1
+ vccd1 _20455_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23173_ _23173_/A vssd1 vssd1 vccd1 vccd1 _27125_/D sky130_fd_sc_hd__clkbuf_1
X_20385_ _20385_/A vssd1 vssd1 vccd1 vccd1 _20385_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22124_ _22124_/A vssd1 vssd1 vccd1 vccd1 _22124_/X sky130_fd_sc_hd__clkbuf_1
X_27981_ _27981_/A _15903_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
XFILLER_122_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22055_ _22071_/A vssd1 vssd1 vccd1 vccd1 _22055_/X sky130_fd_sc_hd__clkbuf_2
X_26932_ _22572_/X _26932_/D vssd1 vssd1 vccd1 vccd1 _26932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21006_ _21006_/A vssd1 vssd1 vccd1 vccd1 _21006_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26863_ _22328_/X _26863_/D vssd1 vssd1 vccd1 vccd1 _26863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25814_ _26013_/CLK _25814_/D vssd1 vssd1 vccd1 vccd1 _25814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26794_ _22082_/X _26794_/D vssd1 vssd1 vccd1 vccd1 _26794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25745_ _25745_/A vssd1 vssd1 vccd1 vccd1 _27829_/D sky130_fd_sc_hd__clkbuf_1
X_22957_ _22957_/A vssd1 vssd1 vccd1 vccd1 _22957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21908_ _21908_/A vssd1 vssd1 vccd1 vccd1 _21908_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13690_ _26901_/Q _13682_/X _13676_/X _13689_/Y vssd1 vssd1 vccd1 vccd1 _26901_/D
+ sky130_fd_sc_hd__a31o_1
X_25676_ _25724_/A vssd1 vssd1 vccd1 vccd1 _25676_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22888_ _22955_/A vssd1 vssd1 vccd1 vccd1 _22888_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27415_ _27415_/CLK _27415_/D vssd1 vssd1 vccd1 vccd1 _27415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24627_ _24627_/A vssd1 vssd1 vccd1 vccd1 _24638_/B sky130_fd_sc_hd__inv_2
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21839_ _21825_/X _21826_/X _21827_/X _21828_/X _21830_/X _21832_/X vssd1 vssd1 vccd1
+ vccd1 _21840_/A sky130_fd_sc_hd__mux4_1
XFILLER_54_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ _14743_/X _26287_/Q _15368_/S vssd1 vssd1 vccd1 vccd1 _15361_/A sky130_fd_sc_hd__mux2_1
X_27346_ _27352_/CLK _27346_/D vssd1 vssd1 vccd1 vccd1 _27346_/Q sky130_fd_sc_hd__dfxtp_2
X_24558_ _24558_/A vssd1 vssd1 vccd1 vccd1 _27540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ _14311_/A vssd1 vssd1 vccd1 vccd1 _14311_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23509_ _23623_/S vssd1 vssd1 vccd1 vccd1 _23525_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_168_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15291_ _26317_/Q _13360_/X _15295_/S vssd1 vssd1 vccd1 vccd1 _15292_/A sky130_fd_sc_hd__mux2_1
X_27277_ _27408_/CLK _27277_/D vssd1 vssd1 vccd1 vccd1 _27277_/Q sky130_fd_sc_hd__dfxtp_1
X_24489_ _24493_/B vssd1 vssd1 vccd1 vccd1 _24505_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ _25914_/Q _25980_/Q _17071_/S vssd1 vssd1 vccd1 vccd1 _17031_/B sky130_fd_sc_hd__mux2_1
X_14242_ _14325_/B vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26228_ _20111_/X _26228_/D vssd1 vssd1 vccd1 vccd1 _26228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14173_ _14225_/A vssd1 vssd1 vccd1 vccd1 _14173_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26159_ _19865_/X _26159_/D vssd1 vssd1 vccd1 vccd1 _26159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13124_ _13124_/A vssd1 vssd1 vccd1 vccd1 _27054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18981_ _18954_/X _18980_/X _18958_/X vssd1 vssd1 vccd1 vccd1 _18981_/X sky130_fd_sc_hd__o21a_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17932_ _18412_/A vssd1 vssd1 vccd1 vccd1 _17932_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13055_ _13142_/B vssd1 vssd1 vccd1 vccd1 _13109_/B sky130_fd_sc_hd__clkbuf_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater108 _27124_/CLK vssd1 vssd1 vccd1 vccd1 _27092_/CLK sky130_fd_sc_hd__clkbuf_1
X_17863_ _18085_/A vssd1 vssd1 vccd1 vccd1 _17863_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater119 _27678_/CLK vssd1 vssd1 vccd1 vccd1 _27285_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19602_ _19602_/A vssd1 vssd1 vccd1 vccd1 _19602_/X sky130_fd_sc_hd__clkbuf_1
X_16814_ _16151_/A _16259_/Y _16260_/X _16261_/X vssd1 vssd1 vccd1 vccd1 _16815_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17794_ _17924_/A vssd1 vssd1 vccd1 vccd1 _18395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_1054 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19533_ _26840_/Q _26808_/Q _26776_/Q _26744_/Q _18788_/X _18790_/X vssd1 vssd1 vccd1
+ vccd1 _19534_/B sky130_fd_sc_hd__mux4_1
X_16745_ _16745_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16765_/B sky130_fd_sc_hd__xnor2_1
X_13957_ _13964_/A vssd1 vssd1 vccd1 vccd1 _14032_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19464_ _19351_/X _19463_/X _19354_/X vssd1 vssd1 vccd1 vccd1 _19464_/X sky130_fd_sc_hd__o21a_1
X_16676_ _16394_/X _16395_/Y _16396_/X vssd1 vssd1 vccd1 vccd1 _16737_/C sky130_fd_sc_hd__a21o_1
X_13888_ _26831_/Q _13880_/X _13886_/X _13887_/Y vssd1 vssd1 vccd1 vccd1 _26831_/D
+ sky130_fd_sc_hd__a31o_1
X_18415_ _18415_/A _18322_/X vssd1 vssd1 vccd1 vccd1 _18415_/X sky130_fd_sc_hd__or2b_1
X_15627_ _15627_/A vssd1 vssd1 vccd1 vccd1 _26169_/D sky130_fd_sc_hd__clkbuf_1
X_19395_ _26161_/Q _26097_/Q _27025_/Q _26993_/Q _19326_/X _19348_/X vssd1 vssd1 vccd1
+ vccd1 _19396_/B sky130_fd_sc_hd__mux4_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18346_ _26286_/Q _26254_/Q _26222_/Q _26190_/Q _18345_/X _18380_/A vssd1 vssd1 vccd1
+ vccd1 _18346_/X sky130_fd_sc_hd__mux4_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _26199_/Q _14718_/A _15562_/S vssd1 vssd1 vccd1 vccd1 _15559_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14509_ _26625_/Q _14496_/X _14492_/X _14508_/Y vssd1 vssd1 vccd1 vccd1 _26625_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18277_ _26155_/Q _26091_/Q _27019_/Q _26987_/Q _18182_/X _18228_/X vssd1 vssd1 vccd1
+ vccd1 _18278_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15489_ _15489_/A vssd1 vssd1 vccd1 vccd1 _26230_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17228_ _25930_/Q _25996_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17229_/B sky130_fd_sc_hd__mux2_1
Xinput30 la1_data_in[29] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_6
Xinput41 la1_oenb[0] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_6
Xinput52 la1_oenb[1] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_4
Xinput63 la1_oenb[2] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17159_ _17220_/A vssd1 vssd1 vccd1 vccd1 _17159_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 wb_clk_i vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_2
XFILLER_157_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20170_ _20162_/X _20163_/X _20164_/X _20165_/X _20167_/X _20169_/X vssd1 vssd1 vccd1
+ vccd1 _20171_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1079 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23860_ _23860_/A vssd1 vssd1 vccd1 vccd1 _23860_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22811_ _22802_/X _22804_/X _22806_/X _22808_/X _22809_/X _22810_/X vssd1 vssd1 vccd1
+ vccd1 _22812_/A sky130_fd_sc_hd__mux4_1
XFILLER_38_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23791_ _27069_/Q _23761_/X _23763_/X _27101_/Q _23765_/X vssd1 vssd1 vccd1 vccd1
+ _23791_/X sky130_fd_sc_hd__a221o_1
XFILLER_16_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25530_ _25560_/A vssd1 vssd1 vccd1 vccd1 _25530_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22742_ _22742_/A vssd1 vssd1 vccd1 vccd1 _22742_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25461_ _25552_/A vssd1 vssd1 vccd1 vccd1 _25461_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22673_ _22665_/X _22666_/X _22667_/X _22668_/X _22669_/X _22670_/X vssd1 vssd1 vccd1
+ vccd1 _22674_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27200_ _27450_/CLK _27200_/D vssd1 vssd1 vccd1 vccd1 _27200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24412_ _24412_/A vssd1 vssd1 vccd1 vccd1 _27485_/D sky130_fd_sc_hd__clkbuf_1
X_21624_ _21624_/A vssd1 vssd1 vccd1 vccd1 _21624_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25392_ _25392_/A vssd1 vssd1 vccd1 vccd1 _27735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27131_ _27827_/CLK _27131_/D vssd1 vssd1 vccd1 vccd1 _27131_/Q sky130_fd_sc_hd__dfxtp_1
X_24343_ _24343_/A vssd1 vssd1 vccd1 vccd1 _27454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1009 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21555_ _21545_/X _21546_/X _21547_/X _21548_/X _21549_/X _21550_/X vssd1 vssd1 vccd1
+ vccd1 _21556_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20506_ _20496_/X _20497_/X _20498_/X _20499_/X _20500_/X _20501_/X vssd1 vssd1 vccd1
+ vccd1 _20507_/A sky130_fd_sc_hd__mux4_1
X_27062_ _23020_/X _27062_/D vssd1 vssd1 vccd1 vccd1 _27062_/Q sky130_fd_sc_hd__dfxtp_1
X_21486_ _21486_/A vssd1 vssd1 vccd1 vccd1 _21486_/X sky130_fd_sc_hd__clkbuf_1
X_24274_ _16194_/X _16196_/Y _16197_/X _24273_/X vssd1 vssd1 vccd1 vccd1 _27411_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26013_ _26013_/CLK _26013_/D vssd1 vssd1 vccd1 vccd1 _26013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23225_ _23225_/A vssd1 vssd1 vccd1 vccd1 _27148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ _20437_/A vssd1 vssd1 vccd1 vccd1 _20437_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23156_ _23167_/A vssd1 vssd1 vccd1 vccd1 _23165_/S sky130_fd_sc_hd__clkbuf_2
X_20368_ _20354_/X _20357_/X _20360_/X _20363_/X _20364_/X _20365_/X vssd1 vssd1 vccd1
+ vccd1 _20369_/A sky130_fd_sc_hd__mux4_1
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22107_ _22543_/A vssd1 vssd1 vccd1 vccd1 _22455_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_23087_ _23087_/A vssd1 vssd1 vccd1 vccd1 _27087_/D sky130_fd_sc_hd__clkbuf_1
X_27964_ _27964_/A _15912_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20299_ _20299_/A vssd1 vssd1 vccd1 vccd1 _20299_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22038_ _22086_/A vssd1 vssd1 vccd1 vccd1 _22038_/X sky130_fd_sc_hd__clkbuf_1
X_26915_ _22510_/X _26915_/D vssd1 vssd1 vccd1 vccd1 _26915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26846_ _22272_/X _26846_/D vssd1 vssd1 vccd1 vccd1 _26846_/Q sky130_fd_sc_hd__dfxtp_1
X_14860_ _26501_/Q _13385_/X _14868_/S vssd1 vssd1 vccd1 vccd1 _14861_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ _26857_/Q _13806_/X _13807_/X _13810_/Y vssd1 vssd1 vccd1 vccd1 _26857_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26777_ _22030_/X _26777_/D vssd1 vssd1 vccd1 vccd1 _26777_/Q sky130_fd_sc_hd__dfxtp_1
X_14791_ _14791_/A vssd1 vssd1 vccd1 vccd1 _14791_/X sky130_fd_sc_hd__clkbuf_2
X_23989_ _23943_/X _23987_/X _23988_/X _23958_/X vssd1 vssd1 vccd1 vccd1 _27295_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16530_ _16289_/A _16400_/A _16067_/X _16528_/Y _16529_/Y vssd1 vssd1 vccd1 vccd1
+ _16623_/C sky130_fd_sc_hd__o221a_1
X_13742_ _26882_/Q _13737_/X _13732_/X _13741_/Y vssd1 vssd1 vccd1 vccd1 _26882_/D
+ sky130_fd_sc_hd__a31o_1
X_25728_ _25728_/A vssd1 vssd1 vccd1 vccd1 _25728_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _16446_/Y _16447_/Y _16460_/Y _25910_/Q vssd1 vssd1 vccd1 vccd1 _16462_/B
+ sky130_fd_sc_hd__a31o_1
X_25659_ _25659_/A vssd1 vssd1 vccd1 vccd1 _25724_/A sky130_fd_sc_hd__clkbuf_2
X_13673_ _15783_/B vssd1 vssd1 vccd1 vccd1 _15190_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18200_ _26824_/Q _26792_/Q _26760_/Q _26728_/Q _18175_/X _18199_/X vssd1 vssd1 vccd1
+ vccd1 _18200_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ _26264_/Q _13325_/X _15418_/S vssd1 vssd1 vccd1 vccd1 _15413_/A sky130_fd_sc_hd__mux2_1
X_19180_ _26696_/Q _26664_/Q _26632_/Q _26600_/Q _19179_/X _19087_/X vssd1 vssd1 vccd1
+ vccd1 _19180_/X sky130_fd_sc_hd__mux4_2
X_16392_ _16674_/A _16715_/B _16715_/C _16737_/B vssd1 vssd1 vccd1 vccd1 _16392_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_730 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18131_ _18127_/X _18130_/X _18197_/S vssd1 vssd1 vccd1 vccd1 _18131_/X sky130_fd_sc_hd__mux2_1
X_27329_ _27402_/CLK _27329_/D vssd1 vssd1 vccd1 vccd1 _27329_/Q sky130_fd_sc_hd__dfxtp_1
X_15343_ _15343_/A vssd1 vssd1 vccd1 vccd1 _26295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18062_ _18384_/A vssd1 vssd1 vccd1 vccd1 _18062_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15274_ _15274_/A vssd1 vssd1 vccd1 vccd1 _26325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17013_ _17013_/A vssd1 vssd1 vccd1 vccd1 _27916_/A sky130_fd_sc_hd__clkbuf_1
X_14225_ _14225_/A vssd1 vssd1 vccd1 vccd1 _14225_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14156_ _26744_/Q _14142_/X _14151_/X _14155_/Y vssd1 vssd1 vccd1 vccd1 _26744_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ _13107_/A vssd1 vssd1 vccd1 vccd1 _27057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14127_/A vssd1 vssd1 vccd1 vccd1 _14098_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ _18952_/X _18959_/X _18963_/X _18866_/X _18840_/X vssd1 vssd1 vccd1 vccd1
+ _18965_/C sky130_fd_sc_hd__a221o_1
XFILLER_98_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17915_ _18014_/A vssd1 vssd1 vccd1 vccd1 _17915_/X sky130_fd_sc_hd__clkbuf_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _14709_/A vssd1 vssd1 vccd1 vccd1 _13038_/X sky130_fd_sc_hd__buf_2
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ _18895_/A vssd1 vssd1 vccd1 vccd1 _18895_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17846_ _18305_/A vssd1 vssd1 vccd1 vccd1 _17846_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17777_ _17777_/A vssd1 vssd1 vccd1 vccd1 _25943_/D sky130_fd_sc_hd__clkbuf_1
X_14989_ _15029_/A vssd1 vssd1 vccd1 vccd1 _14989_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19516_ _19534_/A _19516_/B vssd1 vssd1 vccd1 vccd1 _19516_/X sky130_fd_sc_hd__or2_1
X_16728_ _16728_/A _16780_/B vssd1 vssd1 vccd1 vccd1 _16728_/X sky130_fd_sc_hd__or2_1
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16659_ _16658_/A _16824_/B _16621_/A vssd1 vssd1 vccd1 vccd1 _16659_/Y sky130_fd_sc_hd__o21bai_1
X_19447_ _19444_/X _19446_/X _19468_/S vssd1 vssd1 vccd1 vccd1 _19447_/X sky130_fd_sc_hd__mux2_2
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19378_ _26288_/Q _26256_/Q _26224_/Q _26192_/Q _18778_/X _18782_/X vssd1 vssd1 vccd1
+ vccd1 _19378_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18329_ _18486_/A vssd1 vssd1 vccd1 vccd1 _18329_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21340_ _21340_/A vssd1 vssd1 vccd1 vccd1 _21340_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21271_ _21303_/A vssd1 vssd1 vccd1 vccd1 _21271_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20222_ _20216_/X _20217_/X _20218_/X _20219_/X _20220_/X _20221_/X vssd1 vssd1 vccd1
+ vccd1 _20223_/A sky130_fd_sc_hd__mux4_1
X_23010_ _25636_/A vssd1 vssd1 vccd1 vccd1 _23010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20153_ _20153_/A vssd1 vssd1 vccd1 vccd1 _20153_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20084_ _20076_/X _20077_/X _20078_/X _20079_/X _20081_/X _20083_/X vssd1 vssd1 vccd1
+ vccd1 _20085_/A sky130_fd_sc_hd__mux4_1
X_24961_ _24965_/B _24961_/B vssd1 vssd1 vccd1 vccd1 _24962_/B sky130_fd_sc_hd__or2_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26700_ _21768_/X _26700_/D vssd1 vssd1 vccd1 vccd1 _26700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23912_ _23896_/X _23906_/X _23910_/X _23911_/X vssd1 vssd1 vccd1 vccd1 _27286_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27680_ _27682_/CLK _27680_/D vssd1 vssd1 vccd1 vccd1 _27971_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24892_ _24940_/A vssd1 vssd1 vccd1 vccd1 _24913_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26631_ _21522_/X _26631_/D vssd1 vssd1 vccd1 vccd1 _26631_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23843_ _25921_/Q _25987_/Q _25820_/Q _26019_/Q _23804_/X _23835_/X vssd1 vssd1 vccd1
+ vccd1 _23843_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27949__435 vssd1 vssd1 vccd1 vccd1 _27949__435/HI _27949_/A sky130_fd_sc_hd__conb_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26562_ _21280_/X _26562_/D vssd1 vssd1 vccd1 vccd1 _26562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23774_ _23772_/X _23773_/X _23797_/S vssd1 vssd1 vccd1 vccd1 _23774_/X sky130_fd_sc_hd__mux2_1
X_20986_ _20986_/A vssd1 vssd1 vccd1 vccd1 _20986_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25513_ _25543_/A vssd1 vssd1 vccd1 vccd1 _25513_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22725_ _22716_/X _22718_/X _22720_/X _22722_/X _22723_/X _22724_/X vssd1 vssd1 vccd1
+ vccd1 _22726_/A sky130_fd_sc_hd__mux4_1
XFILLER_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26493_ _21036_/X _26493_/D vssd1 vssd1 vccd1 vccd1 _26493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25444_ _25438_/X _25123_/B _25443_/X _18591_/X vssd1 vssd1 vccd1 vccd1 _25444_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22656_ _22656_/A vssd1 vssd1 vccd1 vccd1 _22656_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21607_ _21599_/X _21600_/X _21601_/X _21602_/X _21603_/X _21604_/X vssd1 vssd1 vccd1
+ vccd1 _21608_/A sky130_fd_sc_hd__mux4_1
X_25375_ _25375_/A vssd1 vssd1 vccd1 vccd1 _27727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22587_ _22577_/X _22578_/X _22579_/X _22580_/X _22581_/X _22582_/X vssd1 vssd1 vccd1
+ vccd1 _22588_/A sky130_fd_sc_hd__mux4_1
XFILLER_182_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27114_ _27127_/CLK _27114_/D vssd1 vssd1 vccd1 vccd1 _27114_/Q sky130_fd_sc_hd__dfxtp_1
X_24326_ _27547_/Q _24328_/B vssd1 vssd1 vccd1 vccd1 _24327_/A sky130_fd_sc_hd__and2_1
X_21538_ _21538_/A vssd1 vssd1 vccd1 vccd1 _21538_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27045_ _22964_/X _27045_/D vssd1 vssd1 vccd1 vccd1 _27045_/Q sky130_fd_sc_hd__dfxtp_1
X_24257_ _24304_/A vssd1 vssd1 vccd1 vccd1 _24264_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_21469_ _21459_/X _21460_/X _21461_/X _21462_/X _21463_/X _21464_/X vssd1 vssd1 vccd1
+ vccd1 _21470_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _14376_/A _14010_/B vssd1 vssd1 vccd1 vccd1 _14010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23208_ _23208_/A vssd1 vssd1 vccd1 vccd1 _27140_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24188_ _24188_/A vssd1 vssd1 vccd1 vccd1 _27364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23139_ _27110_/Q _17715_/X _23143_/S vssd1 vssd1 vccd1 vccd1 _23140_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15961_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15961_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27947_ _27947_/A _15928_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
XFILLER_1_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14912_ _14747_/X _26478_/Q _14918_/S vssd1 vssd1 vccd1 vccd1 _14913_/A sky130_fd_sc_hd__mux2_1
X_17700_ _25919_/Q _17699_/X _17706_/S vssd1 vssd1 vccd1 vccd1 _17701_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18680_ _18680_/A vssd1 vssd1 vccd1 vccd1 _26004_/D sky130_fd_sc_hd__clkbuf_1
X_15892_ _15893_/A vssd1 vssd1 vccd1 vccd1 _15892_/Y sky130_fd_sc_hd__inv_2
X_17631_ _17631_/A vssd1 vssd1 vccd1 vccd1 _25887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14843_ _14843_/A vssd1 vssd1 vccd1 vccd1 _26509_/D sky130_fd_sc_hd__clkbuf_1
X_26829_ _22212_/X _26829_/D vssd1 vssd1 vccd1 vccd1 _26829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ _17469_/X _25857_/Q _17562_/S vssd1 vssd1 vccd1 vccd1 _17563_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ _14774_/A vssd1 vssd1 vccd1 vccd1 _26534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16513_ _16816_/B _16629_/B vssd1 vssd1 vccd1 vccd1 _16664_/A sky130_fd_sc_hd__xnor2_2
X_19301_ _18929_/A _19300_/X _18932_/A vssd1 vssd1 vccd1 vccd1 _19301_/X sky130_fd_sc_hd__o21a_1
XFILLER_189_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13725_ _13904_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13725_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17493_ _17492_/X _25832_/Q _17502_/S vssd1 vssd1 vccd1 vccd1 _17494_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19232_ _27809_/Q _26570_/Q _26442_/Q _26122_/Q _19118_/X _19183_/X vssd1 vssd1 vccd1
+ vccd1 _19232_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16444_ _16780_/B vssd1 vssd1 vccd1 vccd1 _16450_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13656_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19163_ _19161_/X _19162_/X _19211_/S vssd1 vssd1 vccd1 vccd1 _19163_/X sky130_fd_sc_hd__mux2_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _25951_/Q _16375_/B vssd1 vssd1 vccd1 vccd1 _16375_/Y sky130_fd_sc_hd__nand2_1
X_13587_ _13670_/B vssd1 vssd1 vccd1 vccd1 _13587_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18114_ _18114_/A _18066_/X vssd1 vssd1 vccd1 vccd1 _18114_/X sky130_fd_sc_hd__or2b_1
X_15326_ _26301_/Q _13411_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15327_/A sky130_fd_sc_hd__mux2_1
X_19094_ _19091_/X _19092_/X _19211_/S vssd1 vssd1 vccd1 vccd1 _19094_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_28000__466 vssd1 vssd1 vccd1 vccd1 _28000__466/HI _28000_/A sky130_fd_sc_hd__conb_1
X_18045_ _26273_/Q _26241_/Q _26209_/Q _26177_/Q _18044_/X _17937_/X vssd1 vssd1 vccd1
+ vccd1 _18045_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15257_ _15257_/A vssd1 vssd1 vccd1 vccd1 _26332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _14386_/A _14213_/B vssd1 vssd1 vccd1 vccd1 _14208_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15188_ _26362_/Q _13420_/X _15188_/S vssd1 vssd1 vccd1 vccd1 _15189_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ _26750_/Q _14130_/X _14133_/X _14138_/Y vssd1 vssd1 vccd1 vccd1 _26750_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ _20340_/A vssd1 vssd1 vccd1 vccd1 _20065_/A sky130_fd_sc_hd__buf_2
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18947_ _18943_/X _18944_/X _19047_/S vssd1 vssd1 vccd1 vccd1 _18947_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18878_ _18876_/X _18877_/X _19560_/A vssd1 vssd1 vccd1 vccd1 _18878_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17829_ _17924_/A vssd1 vssd1 vccd1 vccd1 _18020_/A sky130_fd_sc_hd__clkbuf_2
X_20840_ _20832_/X _20833_/X _20834_/X _20835_/X _20836_/X _20837_/X vssd1 vssd1 vccd1
+ vccd1 _20841_/A sky130_fd_sc_hd__mux4_1
XFILLER_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20771_ _20771_/A vssd1 vssd1 vccd1 vccd1 _20771_/X sky130_fd_sc_hd__clkbuf_1
X_22510_ _22510_/A vssd1 vssd1 vccd1 vccd1 _22510_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23490_ input27/X _23482_/X _23489_/X _23487_/X vssd1 vssd1 vccd1 vccd1 _27188_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22441_ _22433_/X _22434_/X _22435_/X _22436_/X _22438_/X _22440_/X vssd1 vssd1 vccd1
+ vccd1 _22442_/A sky130_fd_sc_hd__mux4_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1104 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25160_ _27526_/Q _27494_/Q vssd1 vssd1 vccd1 vccd1 _25162_/A sky130_fd_sc_hd__nand2_1
X_22372_ _22436_/A vssd1 vssd1 vccd1 vccd1 _22372_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24111_ _27403_/Q _24117_/B vssd1 vssd1 vccd1 vccd1 _24112_/A sky130_fd_sc_hd__and2_1
XFILLER_159_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21323_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21390_/A sky130_fd_sc_hd__clkbuf_2
X_25091_ _25091_/A vssd1 vssd1 vccd1 vccd1 _27685_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21254_ _21302_/A vssd1 vssd1 vccd1 vccd1 _21254_/X sky130_fd_sc_hd__clkbuf_1
X_24042_ _23849_/A _24040_/X _24041_/X _23864_/A vssd1 vssd1 vccd1 vccd1 _27301_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_606 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20205_ _20237_/A vssd1 vssd1 vccd1 vccd1 _20205_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21185_ _21179_/X _21180_/X _21181_/X _21182_/X _21183_/X _21184_/X vssd1 vssd1 vccd1
+ vccd1 _21186_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27801_ _25652_/X _27801_/D vssd1 vssd1 vccd1 vccd1 _27801_/Q sky130_fd_sc_hd__dfxtp_1
X_20136_ _20130_/X _20131_/X _20132_/X _20133_/X _20134_/X _20135_/X vssd1 vssd1 vccd1
+ vccd1 _20137_/A sky130_fd_sc_hd__mux4_1
XFILLER_131_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25993_ _27145_/CLK _25993_/D vssd1 vssd1 vccd1 vccd1 _25993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27732_ _27746_/CLK _27732_/D vssd1 vssd1 vccd1 vccd1 _27732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20067_ _20067_/A vssd1 vssd1 vccd1 vccd1 _20067_/X sky130_fd_sc_hd__clkbuf_1
X_24944_ _24962_/A _24944_/B vssd1 vssd1 vccd1 vccd1 _24944_/Y sky130_fd_sc_hd__nand2_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27663_ _27663_/CLK _27663_/D vssd1 vssd1 vccd1 vccd1 _27663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24875_ _24889_/A _24875_/B vssd1 vssd1 vccd1 vccd1 _24875_/Y sky130_fd_sc_hd__nand2_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater280 _27592_/CLK vssd1 vssd1 vccd1 vccd1 _27531_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26614_ _21458_/X _26614_/D vssd1 vssd1 vccd1 vccd1 _26614_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater291 _27461_/CLK vssd1 vssd1 vccd1 vccd1 _27562_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23826_ _24014_/A vssd1 vssd1 vccd1 vccd1 _23826_/X sky130_fd_sc_hd__buf_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 _27360_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27594_ _27597_/CLK _27594_/D vssd1 vssd1 vccd1 vccd1 _27594_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_314 _18562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 _21378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_336 _13172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 _13417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26545_ _21220_/X _26545_/D vssd1 vssd1 vccd1 vccd1 _26545_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23757_ _27788_/Q vssd1 vssd1 vccd1 vccd1 _24047_/S sky130_fd_sc_hd__buf_2
XANTENNA_358 _14782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _20953_/X _20954_/X _20955_/X _20956_/X _20958_/X _20960_/X vssd1 vssd1 vccd1
+ vccd1 _20970_/A sky130_fd_sc_hd__mux4_1
XANTENNA_369 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13510_ _13558_/A vssd1 vssd1 vccd1 vccd1 _13510_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22708_ _22708_/A vssd1 vssd1 vccd1 vccd1 _22708_/X sky130_fd_sc_hd__clkbuf_1
X_14490_ _15751_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _14490_/Y sky130_fd_sc_hd__nor2_1
X_26476_ _20984_/X _26476_/D vssd1 vssd1 vccd1 vccd1 _26476_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23688_ _27769_/Q _27249_/Q _23694_/S vssd1 vssd1 vccd1 vccd1 _23689_/A sky130_fd_sc_hd__mux2_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13441_ _14425_/A vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__clkbuf_2
X_25427_ _25427_/A vssd1 vssd1 vccd1 vccd1 _27751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22639_ _22630_/X _22632_/X _22634_/X _22636_/X _22637_/X _22638_/X vssd1 vssd1 vccd1
+ vccd1 _22640_/A sky130_fd_sc_hd__mux4_1
XFILLER_16_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16160_ _16233_/B vssd1 vssd1 vccd1 vccd1 _16249_/B sky130_fd_sc_hd__clkbuf_1
X_13372_ _13372_/A vssd1 vssd1 vccd1 vccd1 _26986_/D sky130_fd_sc_hd__clkbuf_1
X_25358_ _25358_/A _25358_/B vssd1 vssd1 vccd1 vccd1 _25415_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15111_ _15111_/A vssd1 vssd1 vccd1 vccd1 _26397_/D sky130_fd_sc_hd__clkbuf_1
X_24309_ _24309_/A _24384_/B vssd1 vssd1 vccd1 vccd1 _27438_/D sky130_fd_sc_hd__nor2_1
XFILLER_126_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16091_ _16091_/A vssd1 vssd1 vccd1 vccd1 _16738_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25289_ _25273_/A _25282_/A _25288_/X vssd1 vssd1 vccd1 vccd1 _25290_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15042_ _26427_/Q _15040_/X _14966_/B _15041_/Y vssd1 vssd1 vccd1 vccd1 _26427_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27028_ _22904_/X _27028_/D vssd1 vssd1 vccd1 vccd1 _27028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_466 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19850_ _19898_/A vssd1 vssd1 vccd1 vccd1 _19850_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18801_ _19324_/A vssd1 vssd1 vccd1 vccd1 _18801_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19781_ _19813_/A vssd1 vssd1 vccd1 vccd1 _19781_/X sky130_fd_sc_hd__clkbuf_1
X_16993_ input35/X vssd1 vssd1 vccd1 vccd1 _17325_/A sky130_fd_sc_hd__clkbuf_2
X_18732_ _18732_/A vssd1 vssd1 vccd1 vccd1 _26027_/D sky130_fd_sc_hd__clkbuf_1
X_15944_ _15956_/A vssd1 vssd1 vccd1 vccd1 _15949_/A sky130_fd_sc_hd__buf_2
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18663_ _25997_/Q _17737_/X _18663_/S vssd1 vssd1 vccd1 vccd1 _18664_/A sky130_fd_sc_hd__mux2_1
X_15875_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15875_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17614_ _17671_/S vssd1 vssd1 vccd1 vccd1 _17623_/S sky130_fd_sc_hd__clkbuf_2
X_14826_ _14883_/S vssd1 vssd1 vccd1 vccd1 _14835_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_184_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18594_ _18594_/A vssd1 vssd1 vccd1 vccd1 _18594_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ _14756_/X _26539_/Q _14757_/S vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__mux2_1
X_17545_ _17444_/X _25849_/Q _17551_/S vssd1 vssd1 vccd1 vccd1 _17546_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13708_ _13889_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13708_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17476_ _27424_/Q vssd1 vssd1 vccd1 vccd1 _17476_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14688_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14699_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19215_ _19213_/X _19214_/X _19553_/S vssd1 vssd1 vccd1 vccd1 _19215_/X sky130_fd_sc_hd__mux2_2
X_13639_ _13639_/A vssd1 vssd1 vccd1 vccd1 _13639_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16427_ _14779_/A _16384_/X _16375_/B _25954_/Q _16426_/Y vssd1 vssd1 vccd1 vccd1
+ _16786_/B sky130_fd_sc_hd__a221o_2
XFILLER_158_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19146_ _19073_/X _19145_/X _19076_/X vssd1 vssd1 vccd1 vccd1 _19146_/X sky130_fd_sc_hd__o21a_1
X_16358_ _16358_/A vssd1 vssd1 vccd1 vccd1 _16359_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15309_ _26309_/Q _13385_/X _15317_/S vssd1 vssd1 vccd1 vccd1 _15310_/A sky130_fd_sc_hd__mux2_1
X_16289_ _16289_/A _16298_/B _16298_/C vssd1 vssd1 vccd1 vccd1 _16289_/X sky130_fd_sc_hd__or3_1
XFILLER_121_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19077_ _19073_/X _19075_/X _19076_/X vssd1 vssd1 vccd1 vccd1 _19077_/X sky130_fd_sc_hd__o21a_1
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18028_ _18028_/A _18028_/B _18028_/C vssd1 vssd1 vccd1 vccd1 _18029_/A sky130_fd_sc_hd__and3_1
XFILLER_161_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19979_ _19979_/A vssd1 vssd1 vccd1 vccd1 _19979_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22990_ _22990_/A vssd1 vssd1 vccd1 vccd1 _22990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21941_ _21930_/X _21932_/X _21934_/X _21936_/X _21937_/X _21938_/X vssd1 vssd1 vccd1
+ vccd1 _21942_/A sky130_fd_sc_hd__mux4_1
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24660_ _24700_/A vssd1 vssd1 vccd1 vccd1 _24660_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21872_ _21872_/A vssd1 vssd1 vccd1 vccd1 _21872_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23611_ _27781_/Q vssd1 vssd1 vccd1 vccd1 _25601_/A sky130_fd_sc_hd__buf_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _20823_/A vssd1 vssd1 vccd1 vccd1 _20823_/X sky130_fd_sc_hd__clkbuf_1
X_24591_ _24591_/A vssd1 vssd1 vccd1 vccd1 _27555_/D sky130_fd_sc_hd__clkbuf_1
X_26330_ _20471_/X _26330_/D vssd1 vssd1 vccd1 vccd1 _26330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23542_ _24862_/A _27204_/Q _23542_/S vssd1 vssd1 vccd1 vccd1 _23543_/B sky130_fd_sc_hd__mux2_1
X_20754_ _20770_/A vssd1 vssd1 vccd1 vccd1 _20754_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26261_ _20225_/X _26261_/D vssd1 vssd1 vccd1 vccd1 _26261_/Q sky130_fd_sc_hd__dfxtp_1
X_23473_ _27182_/Q _23483_/B vssd1 vssd1 vccd1 vccd1 _23473_/X sky130_fd_sc_hd__or2_1
X_20685_ _20685_/A vssd1 vssd1 vccd1 vccd1 _20685_/X sky130_fd_sc_hd__clkbuf_1
X_28000_ _28000_/A _15880_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_25212_ _25212_/A _25212_/B vssd1 vssd1 vccd1 vccd1 _25213_/B sky130_fd_sc_hd__xor2_1
X_22424_ _22424_/A vssd1 vssd1 vccd1 vccd1 _22424_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26192_ _19983_/X _26192_/D vssd1 vssd1 vccd1 vccd1 _26192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25143_ _25143_/A vssd1 vssd1 vccd1 vccd1 _25309_/A sky130_fd_sc_hd__clkbuf_2
X_22355_ _22347_/X _22348_/X _22349_/X _22350_/X _22352_/X _22354_/X vssd1 vssd1 vccd1
+ vccd1 _22356_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21306_ _21651_/A vssd1 vssd1 vccd1 vccd1 _21377_/A sky130_fd_sc_hd__buf_2
XFILLER_163_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25074_ _25072_/X _25073_/X _25074_/S vssd1 vssd1 vccd1 vccd1 _25074_/X sky130_fd_sc_hd__mux2_1
X_22286_ _22350_/A vssd1 vssd1 vccd1 vccd1 _22286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27992__458 vssd1 vssd1 vccd1 vccd1 _27992__458/HI _27992_/A sky130_fd_sc_hd__conb_1
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24025_ _27094_/Q _27126_/Q _24032_/S vssd1 vssd1 vccd1 vccd1 _24025_/X sky130_fd_sc_hd__mux2_1
X_21237_ _21303_/A vssd1 vssd1 vccd1 vccd1 _21237_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21168_ _21200_/A vssd1 vssd1 vccd1 vccd1 _21168_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20119_ _20151_/A vssd1 vssd1 vccd1 vccd1 _20119_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13990_ _26798_/Q _13987_/X _13983_/X _13989_/Y vssd1 vssd1 vccd1 vccd1 _26798_/D
+ sky130_fd_sc_hd__a31o_1
X_25976_ _27719_/CLK _25976_/D vssd1 vssd1 vccd1 vccd1 _25976_/Q sky130_fd_sc_hd__dfxtp_1
X_21099_ _21093_/X _21094_/X _21095_/X _21096_/X _21097_/X _21098_/X vssd1 vssd1 vccd1
+ vccd1 _21100_/A sky130_fd_sc_hd__mux4_1
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _12941_/A vssd1 vssd1 vccd1 vccd1 _27824_/D sky130_fd_sc_hd__clkbuf_1
X_27715_ _27768_/CLK _27715_/D vssd1 vssd1 vccd1 vccd1 _27715_/Q sky130_fd_sc_hd__dfxtp_1
X_24927_ _24931_/B _24927_/B vssd1 vssd1 vccd1 vccd1 _24928_/B sky130_fd_sc_hd__or2_1
XFILLER_65_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _15660_/A vssd1 vssd1 vccd1 vccd1 _26154_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_100 _19322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24858_ _24867_/C _24858_/B vssd1 vssd1 vccd1 vccd1 _24859_/B sky130_fd_sc_hd__or2_1
X_27646_ _27669_/CLK _27646_/D vssd1 vssd1 vccd1 vccd1 _27646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _20501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _22546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ _26590_/Q _14602_/X _14605_/X _14610_/Y vssd1 vssd1 vccd1 vccd1 _26590_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _24801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23809_ _27071_/Q _27103_/Q _23845_/S vssd1 vssd1 vccd1 vccd1 _23809_/X sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _16017_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15591_ _26184_/Q _14766_/A _15595_/S vssd1 vssd1 vccd1 vccd1 _15592_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27577_ _27577_/CLK _27577_/D vssd1 vssd1 vccd1 vccd1 _27577_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24789_ _24803_/A vssd1 vssd1 vccd1 vccd1 _24800_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_155 _13325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_166 _13401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _25837_/Q _26036_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17330_/X sky130_fd_sc_hd__mux2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _16289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ _15703_/A _14542_/B vssd1 vssd1 vccd1 vccd1 _14542_/Y sky130_fd_sc_hd__nor2_1
X_26528_ _21160_/X _26528_/D vssd1 vssd1 vccd1 vccd1 _26528_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_188 _16495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _14497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _25358_/B vssd1 vssd1 vccd1 vccd1 _17311_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14473_ _26635_/Q _14460_/X _14455_/X _14472_/Y vssd1 vssd1 vccd1 vccd1 _26635_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26459_ _20920_/X _26459_/D vssd1 vssd1 vccd1 vccd1 _26459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19000_ _27799_/Q _26560_/Q _26432_/Q _26112_/Q _18974_/X _18851_/X vssd1 vssd1 vccd1
+ vccd1 _19000_/X sky130_fd_sc_hd__mux4_2
X_16212_ _16212_/A _16221_/B _16235_/C vssd1 vssd1 vccd1 vccd1 _16212_/X sky130_fd_sc_hd__and3_1
X_13424_ _15334_/C _15334_/B _15045_/B vssd1 vssd1 vccd1 vccd1 _13762_/B sky130_fd_sc_hd__or3b_4
X_17192_ _27841_/Q _27145_/Q _25890_/Q _25858_/Q _17142_/X _17191_/X vssd1 vssd1 vccd1
+ vccd1 _17192_/X sky130_fd_sc_hd__mux4_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16143_ _26066_/Q vssd1 vssd1 vccd1 vccd1 _16143_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13355_ _26991_/Q _13353_/X _13367_/S vssd1 vssd1 vccd1 vccd1 _13356_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16074_ _25909_/Q vssd1 vssd1 vccd1 vccd1 _16625_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ _13286_/A vssd1 vssd1 vccd1 vccd1 _27017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15025_ _26434_/Q _15015_/X _15016_/X _15024_/Y vssd1 vssd1 vccd1 vccd1 _26434_/D
+ sky130_fd_sc_hd__a31o_1
X_19902_ _25725_/A vssd1 vssd1 vccd1 vccd1 _19976_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19833_ _19899_/A vssd1 vssd1 vccd1 vccd1 _19833_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19764_ _19812_/A vssd1 vssd1 vccd1 vccd1 _19764_/X sky130_fd_sc_hd__clkbuf_1
X_16976_ _19313_/A _16976_/B vssd1 vssd1 vccd1 vccd1 _16977_/A sky130_fd_sc_hd__and2_1
X_18715_ _18761_/S vssd1 vssd1 vccd1 vccd1 _18724_/S sky130_fd_sc_hd__clkbuf_2
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_15927_ _15930_/A vssd1 vssd1 vccd1 vccd1 _15927_/Y sky130_fd_sc_hd__inv_2
X_19695_ _19727_/A vssd1 vssd1 vccd1 vccd1 _19695_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18646_ _25989_/Q _17712_/X _18652_/S vssd1 vssd1 vccd1 vccd1 _18647_/A sky130_fd_sc_hd__mux2_1
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _15862_/A vssd1 vssd1 vccd1 vccd1 _15858_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ _14809_/A vssd1 vssd1 vccd1 vccd1 _26523_/D sky130_fd_sc_hd__clkbuf_1
X_18577_ _17886_/S _18576_/X _18483_/X vssd1 vssd1 vccd1 vccd1 _18577_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15789_ _15789_/A vssd1 vssd1 vccd1 vccd1 _26104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17528_ _27379_/Q _25735_/B vssd1 vssd1 vccd1 vccd1 _18691_/B sky130_fd_sc_hd__nand2_1
XFILLER_189_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17459_ _17459_/A vssd1 vssd1 vccd1 vccd1 _25821_/D sky130_fd_sc_hd__clkbuf_1
X_28006__472 vssd1 vssd1 vccd1 vccd1 _28006__472/HI _28006_/A sky130_fd_sc_hd__conb_1
XFILLER_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20470_ _20464_/X _20465_/X _20466_/X _20467_/X _20468_/X _20469_/X vssd1 vssd1 vccd1
+ vccd1 _20471_/A sky130_fd_sc_hd__mux4_1
X_19129_ _19123_/X _19125_/X _19128_/X _19035_/X _19105_/X vssd1 vssd1 vccd1 vccd1
+ _19130_/C sky130_fd_sc_hd__a221o_1
XFILLER_173_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22140_ _22140_/A vssd1 vssd1 vccd1 vccd1 _22140_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22071_ _22071_/A vssd1 vssd1 vccd1 vccd1 _22071_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21022_ _21022_/A vssd1 vssd1 vccd1 vccd1 _21022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25830_ _27126_/CLK _25830_/D vssd1 vssd1 vccd1 vccd1 _25830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25761_ _25761_/A vssd1 vssd1 vccd1 vccd1 _27836_/D sky130_fd_sc_hd__clkbuf_1
X_22973_ _25653_/A vssd1 vssd1 vccd1 vccd1 _25635_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27500_ _27747_/CLK _27500_/D vssd1 vssd1 vccd1 vccd1 _27500_/Q sky130_fd_sc_hd__dfxtp_1
X_24712_ _24407_/A _24700_/X _24711_/X _24703_/X vssd1 vssd1 vccd1 vccd1 _27602_/D
+ sky130_fd_sc_hd__o211a_1
X_21924_ _21924_/A vssd1 vssd1 vccd1 vccd1 _21924_/X sky130_fd_sc_hd__clkbuf_1
X_25692_ _25724_/A vssd1 vssd1 vccd1 vccd1 _25692_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27431_ _27436_/CLK _27431_/D vssd1 vssd1 vccd1 vccd1 _27431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24643_ _24700_/A vssd1 vssd1 vccd1 vccd1 _24643_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21855_ _21844_/X _21846_/X _21848_/X _21850_/X _21851_/X _21852_/X vssd1 vssd1 vccd1
+ vccd1 _21856_/A sky130_fd_sc_hd__mux4_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _20791_/X _20795_/X _20799_/X _20803_/X _20804_/X _20805_/X vssd1 vssd1 vccd1
+ vccd1 _20807_/A sky130_fd_sc_hd__mux4_1
X_27362_ _27825_/CLK _27362_/D vssd1 vssd1 vccd1 vccd1 _27362_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24574_ _27648_/Q _24576_/B vssd1 vssd1 vccd1 vccd1 _24575_/A sky130_fd_sc_hd__and2_1
X_21786_ _21786_/A vssd1 vssd1 vccd1 vccd1 _21786_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26313_ _20405_/X _26313_/D vssd1 vssd1 vccd1 vccd1 _26313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23525_ _24835_/A _27199_/Q _23525_/S vssd1 vssd1 vccd1 vccd1 _23526_/B sky130_fd_sc_hd__mux2_1
X_27293_ _27293_/CLK _27293_/D vssd1 vssd1 vccd1 vccd1 _27293_/Q sky130_fd_sc_hd__dfxtp_1
X_20737_ _20737_/A vssd1 vssd1 vccd1 vccd1 _20737_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26244_ _20161_/X _26244_/D vssd1 vssd1 vccd1 vccd1 _26244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23456_ _27176_/Q _23456_/B vssd1 vssd1 vccd1 vccd1 _23456_/X sky130_fd_sc_hd__or2_1
XFILLER_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20668_ _20684_/A vssd1 vssd1 vccd1 vccd1 _20668_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22407_ _22401_/X _22402_/X _22403_/X _22404_/X _22405_/X _22406_/X vssd1 vssd1 vccd1
+ vccd1 _22408_/A sky130_fd_sc_hd__mux4_1
XFILLER_52_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26175_ _19931_/X _26175_/D vssd1 vssd1 vccd1 vccd1 _26175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23387_ _27779_/Q vssd1 vssd1 vccd1 vccd1 _24804_/A sky130_fd_sc_hd__inv_2
X_20599_ _20599_/A vssd1 vssd1 vccd1 vccd1 _20599_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25126_ _27522_/Q _27490_/Q vssd1 vssd1 vccd1 vccd1 _25126_/X sky130_fd_sc_hd__or2_1
X_13140_ _27051_/Q _13139_/X _13140_/S vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__mux2_1
X_22338_ _22338_/A vssd1 vssd1 vccd1 vccd1 _22338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25057_ _27075_/Q _27107_/Q _25088_/S vssd1 vssd1 vccd1 vccd1 _25057_/X sky130_fd_sc_hd__mux2_1
X_13071_ _27363_/Q _13063_/X _13064_/X _27331_/Q _13070_/X vssd1 vssd1 vccd1 vccd1
+ _14721_/A sky130_fd_sc_hd__a221o_2
X_22269_ _22261_/X _22262_/X _22263_/X _22264_/X _22266_/X _22268_/X vssd1 vssd1 vccd1
+ vccd1 _22270_/A sky130_fd_sc_hd__mux4_1
XFILLER_183_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24008_ _25938_/Q _26004_/Q _25837_/Q _26036_/Q _23993_/X _23976_/X vssd1 vssd1 vccd1
+ vccd1 _24008_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16830_ _16561_/A _16648_/C _16829_/X _16797_/A vssd1 vssd1 vccd1 vccd1 _16830_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_120_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_527 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13973_ _16563_/A vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__buf_2
XFILLER_111_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16761_ _16342_/Y _16761_/B _16862_/A vssd1 vssd1 vccd1 vccd1 _16761_/X sky130_fd_sc_hd__and3b_1
X_25959_ _26056_/CLK _25959_/D vssd1 vssd1 vccd1 vccd1 _25959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18500_ _18468_/X _18495_/X _18499_/X _18412_/X vssd1 vssd1 vccd1 vccd1 _18509_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1186 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15712_ _15712_/A vssd1 vssd1 vccd1 vccd1 _15766_/A sky130_fd_sc_hd__clkbuf_2
X_12924_ input71/X input72/X input42/X input43/X vssd1 vssd1 vccd1 vccd1 _12928_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_74_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19480_ _19478_/X _19479_/X _19480_/S vssd1 vssd1 vccd1 vccd1 _19480_/X sky130_fd_sc_hd__mux2_1
X_16692_ _16692_/A _16692_/B _16692_/C vssd1 vssd1 vccd1 vccd1 _16692_/X sky130_fd_sc_hd__or3_1
X_18431_ _26706_/Q _26674_/Q _26642_/Q _26610_/Q _18360_/X _18408_/X vssd1 vssd1 vccd1
+ vccd1 _18432_/A sky130_fd_sc_hd__mux4_1
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27629_ _27629_/CLK _27629_/D vssd1 vssd1 vccd1 vccd1 _27629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15643_ _13105_/X _26161_/Q _15645_/S vssd1 vssd1 vccd1 vccd1 _15644_/A sky130_fd_sc_hd__mux2_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _18362_/A _18317_/X vssd1 vssd1 vccd1 vccd1 _18362_/X sky130_fd_sc_hd__or2b_1
X_15574_ _15574_/A vssd1 vssd1 vccd1 vccd1 _26192_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17313_ input36/X vssd1 vssd1 vccd1 vccd1 _17313_/X sky130_fd_sc_hd__clkbuf_2
X_14525_ _15777_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14525_/Y sky130_fd_sc_hd__nor2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18293_ _18293_/A _17910_/X vssd1 vssd1 vccd1 vccd1 _18293_/X sky130_fd_sc_hd__or2b_1
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17244_ _17242_/X _17243_/X _17220_/X vssd1 vssd1 vccd1 vccd1 _17244_/X sky130_fd_sc_hd__a21bo_1
X_14456_ _16289_/A vssd1 vssd1 vccd1 vccd1 _15728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13407_ _13407_/A vssd1 vssd1 vccd1 vccd1 _26975_/D sky130_fd_sc_hd__clkbuf_1
X_17175_ _27208_/Q _17174_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17176_/A sky130_fd_sc_hd__mux2_1
X_14387_ _26661_/Q _14379_/X _14385_/X _14386_/Y vssd1 vssd1 vccd1 vccd1 _26661_/D
+ sky130_fd_sc_hd__a31o_1
X_16126_ _26071_/Q vssd1 vssd1 vccd1 vccd1 _16126_/Y sky130_fd_sc_hd__inv_2
X_13338_ _13421_/S vssd1 vssd1 vccd1 vccd1 _13351_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_6_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ _16056_/Y _13425_/A _27266_/Q _16047_/Y vssd1 vssd1 vccd1 vccd1 _16057_/X
+ sky130_fd_sc_hd__a22o_1
X_13269_ _27024_/Q _13111_/X _13269_/S vssd1 vssd1 vccd1 vccd1 _13270_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15008_ _15745_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _15008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19816_ _25725_/A vssd1 vssd1 vccd1 vccd1 _19886_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19747_ _19813_/A vssd1 vssd1 vccd1 vccd1 _19747_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_398 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16959_ _27582_/Q _24636_/B vssd1 vssd1 vccd1 vccd1 _16960_/A sky130_fd_sc_hd__and2_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19678_ _19726_/A vssd1 vssd1 vccd1 vccd1 _19678_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18629_ _18629_/A vssd1 vssd1 vccd1 vccd1 _25981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21640_ _21640_/A vssd1 vssd1 vccd1 vccd1 _21640_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21571_ _21561_/X _21562_/X _21563_/X _21564_/X _21566_/X _21568_/X vssd1 vssd1 vccd1
+ vccd1 _21572_/A sky130_fd_sc_hd__mux4_1
XANTENNA_11 _25856_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_22 _27141_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23310_ _27724_/Q _23290_/Y _27748_/Q _23261_/Y vssd1 vssd1 vccd1 vccd1 _23310_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_33 _17714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20522_ _20512_/X _20513_/X _20514_/X _20515_/X _20517_/X _20519_/X vssd1 vssd1 vccd1
+ vccd1 _20523_/A sky130_fd_sc_hd__mux4_1
XANTENNA_44 _17921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24290_ _24290_/A _24317_/B vssd1 vssd1 vccd1 vccd1 _24291_/A sky130_fd_sc_hd__and2_1
XFILLER_21_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_55 _18218_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_66 _18331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23241_ _23241_/A vssd1 vssd1 vccd1 vccd1 _27155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_77 _18524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_88 _18920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20453_ _20501_/A vssd1 vssd1 vccd1 vccd1 _20453_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_99 _19309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23172_ _27125_/Q _17763_/X _23176_/S vssd1 vssd1 vccd1 vccd1 _23173_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20384_ _20376_/X _20377_/X _20378_/X _20379_/X _20380_/X _20381_/X vssd1 vssd1 vccd1
+ vccd1 _20385_/A sky130_fd_sc_hd__mux4_1
XFILLER_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22123_ _22103_/X _22106_/X _22109_/X _22112_/X _22113_/X _22114_/X vssd1 vssd1 vccd1
+ vccd1 _22124_/A sky130_fd_sc_hd__mux4_1
XFILLER_134_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27980_ _27980_/A _15904_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
XFILLER_88_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22054_ _22086_/A vssd1 vssd1 vccd1 vccd1 _22054_/X sky130_fd_sc_hd__clkbuf_1
X_26931_ _22570_/X _26931_/D vssd1 vssd1 vccd1 vccd1 _26931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21005_ _20991_/X _20992_/X _20993_/X _20994_/X _20995_/X _20996_/X vssd1 vssd1 vccd1
+ vccd1 _21006_/A sky130_fd_sc_hd__mux4_1
XFILLER_47_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26862_ _22326_/X _26862_/D vssd1 vssd1 vccd1 vccd1 _26862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25813_ _26013_/CLK _25813_/D vssd1 vssd1 vccd1 vccd1 _25813_/Q sky130_fd_sc_hd__dfxtp_1
X_26793_ _22080_/X _26793_/D vssd1 vssd1 vccd1 vccd1 _26793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25744_ _17434_/X _27829_/Q _25746_/S vssd1 vssd1 vccd1 vccd1 _25745_/A sky130_fd_sc_hd__mux2_1
X_22956_ _22956_/A vssd1 vssd1 vccd1 vccd1 _22956_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21907_ _21895_/X _21896_/X _21897_/X _21898_/X _21899_/X _21900_/X vssd1 vssd1 vccd1
+ vccd1 _21908_/A sky130_fd_sc_hd__mux4_1
XFILLER_56_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25675_ _25723_/A vssd1 vssd1 vccd1 vccd1 _25675_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22887_ _22887_/A vssd1 vssd1 vccd1 vccd1 _22955_/A sky130_fd_sc_hd__buf_2
XFILLER_102_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24626_ _27584_/Q _27583_/Q _24635_/B _24626_/D vssd1 vssd1 vccd1 vccd1 _24627_/A
+ sky130_fd_sc_hd__or4_1
X_27414_ _27414_/CLK _27414_/D vssd1 vssd1 vccd1 vccd1 _27414_/Q sky130_fd_sc_hd__dfxtp_1
X_21838_ _21838_/A vssd1 vssd1 vccd1 vccd1 _21838_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27345_ _27352_/CLK _27345_/D vssd1 vssd1 vccd1 vccd1 _27345_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24557_ _27640_/Q _24565_/B vssd1 vssd1 vccd1 vccd1 _24558_/A sky130_fd_sc_hd__and2_1
XFILLER_197_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21769_ _21758_/X _21760_/X _21762_/X _21764_/X _21765_/X _21766_/X vssd1 vssd1 vccd1
+ vccd1 _21770_/A sky130_fd_sc_hd__mux4_1
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _14365_/A vssd1 vssd1 vccd1 vccd1 _14310_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23508_ _23600_/A vssd1 vssd1 vccd1 vccd1 _23623_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_196_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15290_ _15290_/A vssd1 vssd1 vccd1 vccd1 _26318_/D sky130_fd_sc_hd__clkbuf_1
X_27276_ _27278_/CLK _27276_/D vssd1 vssd1 vccd1 vccd1 _27276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24488_ _27583_/Q _24488_/B vssd1 vssd1 vccd1 vccd1 _24493_/B sky130_fd_sc_hd__nand2_1
X_27998__464 vssd1 vssd1 vccd1 vccd1 _27998__464/HI _27998_/A sky130_fd_sc_hd__conb_1
X_14241_ _14257_/A vssd1 vssd1 vccd1 vccd1 _14325_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26227_ _20109_/X _26227_/D vssd1 vssd1 vccd1 vccd1 _26227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23439_ _17048_/S _23429_/X _23438_/X _23434_/X vssd1 vssd1 vccd1 vccd1 _27169_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14172_ _14172_/A vssd1 vssd1 vccd1 vccd1 _14225_/A sky130_fd_sc_hd__buf_2
X_26158_ _19863_/X _26158_/D vssd1 vssd1 vccd1 vccd1 _26158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25109_ _25733_/A _18594_/X _27753_/D _25108_/Y vssd1 vssd1 vccd1 vccd1 _27688_/D
+ sky130_fd_sc_hd__o211a_1
X_13123_ _27054_/Q _13122_/X _13140_/S vssd1 vssd1 vccd1 vccd1 _13124_/A sky130_fd_sc_hd__mux2_1
XFILLER_180_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26089_ _19620_/X _26089_/D vssd1 vssd1 vccd1 vccd1 _26089_/Q sky130_fd_sc_hd__dfxtp_1
X_18980_ _26271_/Q _26239_/Q _26207_/Q _26175_/Q _18859_/X _18955_/X vssd1 vssd1 vccd1
+ vccd1 _18980_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _17888_/X _17927_/X _17930_/X _17894_/X vssd1 vssd1 vccd1 vccd1 _17931_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13054_ _13169_/B vssd1 vssd1 vccd1 vccd1 _13142_/B sky130_fd_sc_hd__clkbuf_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17862_ _17860_/X _17861_/X _17886_/S vssd1 vssd1 vccd1 vccd1 _17862_/X sky130_fd_sc_hd__mux2_1
Xrepeater109 _27123_/CLK vssd1 vssd1 vccd1 vccd1 _27124_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_121_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19601_ _19589_/X _19590_/X _19591_/X _19592_/X _19593_/X _19594_/X vssd1 vssd1 vccd1
+ vccd1 _19602_/A sky130_fd_sc_hd__mux4_1
X_16813_ _16777_/X _16782_/X _16788_/X _16844_/A vssd1 vssd1 vccd1 vccd1 _16841_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_495 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17793_ _27595_/Q vssd1 vssd1 vccd1 vccd1 _17924_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_143_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19532_ _19532_/A vssd1 vssd1 vccd1 vccd1 _26071_/D sky130_fd_sc_hd__clkbuf_1
X_16744_ _16744_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16744_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_1040 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13956_ _16134_/A vssd1 vssd1 vccd1 vccd1 _14340_/A sky130_fd_sc_hd__buf_2
XFILLER_93_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19463_ _26292_/Q _26260_/Q _26228_/Q _26196_/Q _19441_/X _19352_/X vssd1 vssd1 vccd1
+ vccd1 _19463_/X sky130_fd_sc_hd__mux4_1
X_13887_ _13887_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13887_/Y sky130_fd_sc_hd__nor2_1
X_16675_ _16852_/A _16715_/B vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__or2_1
XFILLER_62_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18414_ _26161_/Q _26097_/Q _27025_/Q _26993_/Q _18298_/X _18387_/X vssd1 vssd1 vccd1
+ vccd1 _18415_/A sky130_fd_sc_hd__mux4_2
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _13038_/X _26169_/Q _15634_/S vssd1 vssd1 vccd1 vccd1 _15627_/A sky130_fd_sc_hd__mux2_1
X_19394_ _19384_/X _19388_/X _19392_/X _19324_/X _19393_/X vssd1 vssd1 vccd1 vccd1
+ _19405_/B sky130_fd_sc_hd__a221o_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18345_ _18360_/A vssd1 vssd1 vccd1 vccd1 _18345_/X sky130_fd_sc_hd__buf_4
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15557_/A vssd1 vssd1 vccd1 vccd1 _26200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14508_ _15764_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14508_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18276_ _18150_/X _18271_/X _18275_/X _18253_/X vssd1 vssd1 vccd1 vccd1 _18287_/B
+ sky130_fd_sc_hd__a211o_1
X_15488_ _13072_/X _26230_/Q _15490_/S vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 la1_data_in[1] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_4
X_17227_ _27844_/Q _27148_/Q _25893_/Q _25861_/Q _17203_/X _17191_/X vssd1 vssd1 vccd1
+ vccd1 _17227_/X sky130_fd_sc_hd__mux4_1
X_14439_ _15714_/A _14446_/B vssd1 vssd1 vccd1 vccd1 _14439_/Y sky130_fd_sc_hd__nor2_1
Xinput31 la1_data_in[2] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 la1_oenb[10] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_2
Xinput53 la1_oenb[20] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_2
Xinput64 la1_oenb[30] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_4
X_17158_ _25823_/Q _26022_/Q _17158_/S vssd1 vssd1 vccd1 vccd1 _17158_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16109_ _16109_/A vssd1 vssd1 vccd1 vccd1 _16110_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17089_ _27072_/Q _27104_/Q _17112_/S vssd1 vssd1 vccd1 vccd1 _17089_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22810_ _22858_/A vssd1 vssd1 vccd1 vccd1 _22810_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23790_ _23788_/X _23789_/X _23797_/S vssd1 vssd1 vccd1 vccd1 _23790_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22741_ _22735_/X _22736_/X _22737_/X _22738_/X _22739_/X _22740_/X vssd1 vssd1 vccd1
+ vccd1 _22742_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25460_ _27694_/Q _25448_/X _25449_/X vssd1 vssd1 vccd1 vccd1 _25460_/Y sky130_fd_sc_hd__a21oi_1
X_22672_ _22672_/A vssd1 vssd1 vccd1 vccd1 _22672_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24411_ _27586_/Q _24411_/B vssd1 vssd1 vccd1 vccd1 _24412_/A sky130_fd_sc_hd__and2_1
XFILLER_197_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21623_ _21615_/X _21616_/X _21617_/X _21618_/X _21619_/X _21620_/X vssd1 vssd1 vccd1
+ vccd1 _21624_/A sky130_fd_sc_hd__mux4_1
XFILLER_34_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25391_ _27735_/Q input46/X _25391_/S vssd1 vssd1 vccd1 vccd1 _25392_/A sky130_fd_sc_hd__mux2_1
X_27130_ _27130_/CLK _27130_/D vssd1 vssd1 vccd1 vccd1 _27130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24342_ _27554_/Q _24350_/B vssd1 vssd1 vccd1 vccd1 _24343_/A sky130_fd_sc_hd__and2_1
X_21554_ _21554_/A vssd1 vssd1 vccd1 vccd1 _21554_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20505_ _20505_/A vssd1 vssd1 vccd1 vccd1 _20505_/X sky130_fd_sc_hd__clkbuf_1
X_27061_ _23018_/X _27061_/D vssd1 vssd1 vccd1 vccd1 _27061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24273_ _24279_/A vssd1 vssd1 vccd1 vccd1 _24273_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21485_ _21475_/X _21476_/X _21477_/X _21478_/X _21480_/X _21482_/X vssd1 vssd1 vccd1
+ vccd1 _21486_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26012_ _26012_/CLK _26012_/D vssd1 vssd1 vccd1 vccd1 _26012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23224_ _17482_/X _27148_/Q _23226_/S vssd1 vssd1 vccd1 vccd1 _23225_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20436_ _20424_/X _20425_/X _20426_/X _20427_/X _20430_/X _20433_/X vssd1 vssd1 vccd1
+ vccd1 _20437_/A sky130_fd_sc_hd__mux4_1
XFILLER_14_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23155_ _23155_/A vssd1 vssd1 vccd1 vccd1 _27117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20367_ _20367_/A vssd1 vssd1 vccd1 vccd1 _20367_/X sky130_fd_sc_hd__clkbuf_1
X_22106_ _22174_/A vssd1 vssd1 vccd1 vccd1 _22106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23086_ _27087_/Q _17744_/X _23092_/S vssd1 vssd1 vccd1 vccd1 _23087_/A sky130_fd_sc_hd__mux2_1
X_27963_ _27963_/A _15864_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
X_20298_ _20286_/X _20287_/X _20288_/X _20289_/X _20290_/X _20291_/X vssd1 vssd1 vccd1
+ vccd1 _20299_/A sky130_fd_sc_hd__mux4_1
X_22037_ _22085_/A vssd1 vssd1 vccd1 vccd1 _22037_/X sky130_fd_sc_hd__clkbuf_1
X_26914_ _22502_/X _26914_/D vssd1 vssd1 vccd1 vccd1 _26914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26845_ _22270_/X _26845_/D vssd1 vssd1 vccd1 vccd1 _26845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13810_ _13902_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13810_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14790_ _14790_/A vssd1 vssd1 vccd1 vccd1 _26529_/D sky130_fd_sc_hd__clkbuf_1
X_23988_ _27090_/Q _23954_/X _23955_/X _27122_/Q _23956_/X vssd1 vssd1 vccd1 vccd1
+ _23988_/X sky130_fd_sc_hd__a221o_1
X_26776_ _22028_/X _26776_/D vssd1 vssd1 vccd1 vccd1 _26776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ _13921_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13741_/Y sky130_fd_sc_hd__nor2_1
X_25727_ _25721_/X _25722_/X _25723_/X _25724_/X _25725_/X _25726_/X vssd1 vssd1 vccd1
+ vccd1 _25728_/A sky130_fd_sc_hd__mux4_1
X_22939_ _22955_/A vssd1 vssd1 vccd1 vccd1 _22939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ _13672_/A _13672_/B _13425_/A vssd1 vssd1 vccd1 vccd1 _15783_/B sky130_fd_sc_hd__or3b_4
X_16460_ _16728_/A _16460_/B vssd1 vssd1 vccd1 vccd1 _16460_/Y sky130_fd_sc_hd__nor2_1
X_25658_ _25723_/A vssd1 vssd1 vccd1 vccd1 _25658_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15411_ _15411_/A vssd1 vssd1 vccd1 vccd1 _26265_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24609_ _27664_/Q _24609_/B vssd1 vssd1 vccd1 vccd1 _24610_/A sky130_fd_sc_hd__and2_1
X_16391_ _16742_/A _16393_/B vssd1 vssd1 vccd1 vccd1 _16737_/B sky130_fd_sc_hd__xnor2_2
XFILLER_185_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25589_ _25572_/X _25582_/X _25583_/X _24949_/B _25584_/X vssd1 vssd1 vccd1 vccd1
+ _25589_/X sky130_fd_sc_hd__o311a_1
XFILLER_197_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18130_ _26949_/Q _26917_/Q _26885_/Q _26853_/Q _18101_/X _18129_/X vssd1 vssd1 vccd1
+ vccd1 _18130_/X sky130_fd_sc_hd__mux4_2
X_15342_ _14718_/X _26295_/Q _15346_/S vssd1 vssd1 vccd1 vccd1 _15343_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27328_ _27328_/CLK _27328_/D vssd1 vssd1 vccd1 vccd1 _27328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_742 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18061_ _18061_/A _17978_/X vssd1 vssd1 vccd1 vccd1 _18061_/X sky130_fd_sc_hd__or2b_1
X_15273_ _26325_/Q _13334_/X _15273_/S vssd1 vssd1 vccd1 vccd1 _15274_/A sky130_fd_sc_hd__mux2_1
X_27259_ _27261_/CLK _27259_/D vssd1 vssd1 vccd1 vccd1 _27259_/Q sky130_fd_sc_hd__dfxtp_1
X_14224_ _26719_/Q _14212_/X _14220_/X _14223_/Y vssd1 vssd1 vccd1 vccd1 _26719_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17012_ _27195_/Q _17007_/X _17067_/S vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14155_ _14333_/A _14158_/B vssd1 vssd1 vccd1 vccd1 _14155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13106_ _27057_/Q _13105_/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14086_ _26770_/Q _14076_/X _14080_/X _14085_/Y vssd1 vssd1 vccd1 vccd1 _26770_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18963_ _18960_/X _18961_/X _19057_/S vssd1 vssd1 vccd1 vccd1 _18963_/X sky130_fd_sc_hd__mux2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17914_ _26268_/Q _26236_/Q _26204_/Q _26172_/Q _17801_/X _17913_/X vssd1 vssd1 vccd1
+ vccd1 _17914_/X sky130_fd_sc_hd__mux4_2
X_13037_ _27366_/Q _13022_/X _13030_/X _27334_/Q _13036_/X vssd1 vssd1 vccd1 vccd1
+ _14709_/A sky130_fd_sc_hd__a221o_1
XFILLER_152_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18894_ _19448_/A vssd1 vssd1 vccd1 vccd1 _18895_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17845_ _17898_/A vssd1 vssd1 vccd1 vccd1 _18305_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ _25943_/Q _17775_/X _17776_/S vssd1 vssd1 vccd1 vccd1 _17777_/A sky130_fd_sc_hd__mux2_1
X_14988_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14988_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19515_ _26839_/Q _26807_/Q _26775_/Q _26743_/Q _18788_/X _19407_/X vssd1 vssd1 vccd1
+ vccd1 _19516_/B sky130_fd_sc_hd__mux4_1
X_16727_ _16450_/Y _16481_/A _16606_/Y _16641_/A vssd1 vssd1 vccd1 vccd1 _16727_/X
+ sky130_fd_sc_hd__a31o_1
X_13939_ _26811_/Q _13933_/X _13861_/B _13938_/Y vssd1 vssd1 vccd1 vccd1 _26811_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19446_ _26547_/Q _26515_/Q _26483_/Q _27059_/Q _19401_/X _19445_/X vssd1 vssd1 vccd1
+ vccd1 _19446_/X sky130_fd_sc_hd__mux4_1
X_16658_ _16658_/A _16824_/B vssd1 vssd1 vccd1 vccd1 _16658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _26176_/Q _14791_/A _15617_/S vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__mux2_1
X_19377_ _19555_/A _19377_/B vssd1 vssd1 vccd1 vccd1 _19377_/X sky130_fd_sc_hd__or2_1
X_16589_ _16578_/Y _16636_/B _16913_/B vssd1 vssd1 vccd1 vccd1 _16879_/B sky130_fd_sc_hd__o21a_1
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18328_ _26541_/Q _26509_/Q _26477_/Q _27053_/Q _18233_/X _18259_/X vssd1 vssd1 vccd1
+ vccd1 _18328_/X sky130_fd_sc_hd__mux4_1
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18259_ _18418_/A vssd1 vssd1 vccd1 vccd1 _18259_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21270_ _21302_/A vssd1 vssd1 vccd1 vccd1 _21270_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20221_ _20237_/A vssd1 vssd1 vccd1 vccd1 _20221_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20152_ _20146_/X _20147_/X _20148_/X _20149_/X _20150_/X _20151_/X vssd1 vssd1 vccd1
+ vccd1 _20153_/A sky130_fd_sc_hd__mux4_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24960_ _24960_/A _24960_/B vssd1 vssd1 vccd1 vccd1 _24961_/B sky130_fd_sc_hd__nor2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _20151_/A vssd1 vssd1 vccd1 vccd1 _20083_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23911_ _24005_/A vssd1 vssd1 vccd1 vccd1 _23911_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24891_ _27654_/Q _24885_/X _24889_/Y _24890_/X vssd1 vssd1 vccd1 vccd1 _27654_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26630_ _21520_/X _26630_/D vssd1 vssd1 vccd1 vccd1 _26630_/Q sky130_fd_sc_hd__dfxtp_1
X_23842_ _27835_/Q _27139_/Q _25884_/Q _25852_/Q _23826_/X _23802_/X vssd1 vssd1 vccd1
+ vccd1 _23842_/X sky130_fd_sc_hd__mux4_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26561_ _21278_/X _26561_/D vssd1 vssd1 vccd1 vccd1 _26561_/Q sky130_fd_sc_hd__dfxtp_1
X_23773_ _27067_/Q _27099_/Q _23796_/S vssd1 vssd1 vccd1 vccd1 _23773_/X sky130_fd_sc_hd__mux2_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20985_ _20972_/X _20974_/X _20976_/X _20978_/X _20979_/X _20980_/X vssd1 vssd1 vccd1
+ vccd1 _20986_/A sky130_fd_sc_hd__mux4_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25512_ _25487_/X _25492_/X _25493_/X _24883_/B _25494_/X vssd1 vssd1 vccd1 vccd1
+ _25512_/X sky130_fd_sc_hd__o311a_1
XFILLER_53_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22724_ _22772_/A vssd1 vssd1 vccd1 vccd1 _22724_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26492_ _21034_/X _26492_/D vssd1 vssd1 vccd1 vccd1 _26492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25443_ _24267_/A _25440_/X _25442_/X _25524_/A _24831_/B vssd1 vssd1 vccd1 vccd1
+ _25443_/X sky130_fd_sc_hd__o311a_1
X_22655_ _22649_/X _22650_/X _22651_/X _22652_/X _22653_/X _22654_/X vssd1 vssd1 vccd1
+ vccd1 _22656_/A sky130_fd_sc_hd__mux4_1
XFILLER_41_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21606_ _21606_/A vssd1 vssd1 vccd1 vccd1 _21606_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25374_ _27727_/Q input69/X _25380_/S vssd1 vssd1 vccd1 vccd1 _25375_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22586_ _22586_/A vssd1 vssd1 vccd1 vccd1 _22586_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27113_ _27856_/CLK _27113_/D vssd1 vssd1 vccd1 vccd1 _27113_/Q sky130_fd_sc_hd__dfxtp_1
X_24325_ _24325_/A vssd1 vssd1 vccd1 vccd1 _27446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21537_ _21529_/X _21530_/X _21531_/X _21532_/X _21533_/X _21534_/X vssd1 vssd1 vccd1
+ vccd1 _21538_/A sky130_fd_sc_hd__mux4_1
XFILLER_181_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27044_ _22954_/X _27044_/D vssd1 vssd1 vccd1 vccd1 _27044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24256_ _24256_/A _24256_/B vssd1 vssd1 vccd1 vccd1 _27400_/D sky130_fd_sc_hd__nor2_1
XFILLER_107_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21468_ _21468_/A vssd1 vssd1 vccd1 vccd1 _21468_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23207_ _17456_/X _27140_/Q _23215_/S vssd1 vssd1 vccd1 vccd1 _23208_/A sky130_fd_sc_hd__mux2_1
X_20419_ _20419_/A vssd1 vssd1 vccd1 vccd1 _20419_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24187_ _27469_/Q _24195_/B vssd1 vssd1 vccd1 vccd1 _24188_/A sky130_fd_sc_hd__and2_1
X_21399_ _21389_/X _21390_/X _21391_/X _21392_/X _21394_/X _21396_/X vssd1 vssd1 vccd1
+ vccd1 _21400_/A sky130_fd_sc_hd__mux4_1
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23138_ _23138_/A vssd1 vssd1 vccd1 vccd1 _27109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23069_ _23069_/A vssd1 vssd1 vccd1 vccd1 _27079_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27946_ _27946_/A _15929_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
X_15960_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15960_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14911_ _14911_/A vssd1 vssd1 vccd1 vccd1 _26479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15891_ _15893_/A vssd1 vssd1 vccd1 vccd1 _15891_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17630_ _17463_/X _25887_/Q _17634_/S vssd1 vssd1 vccd1 vccd1 _17631_/A sky130_fd_sc_hd__mux2_1
X_26828_ _22210_/X _26828_/D vssd1 vssd1 vccd1 vccd1 _26828_/Q sky130_fd_sc_hd__dfxtp_1
X_14842_ _26509_/Q _13360_/X _14846_/S vssd1 vssd1 vccd1 vccd1 _14843_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17561_ _17561_/A vssd1 vssd1 vccd1 vccd1 _25856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26759_ _21964_/X _26759_/D vssd1 vssd1 vccd1 vccd1 _26759_/Q sky130_fd_sc_hd__dfxtp_1
X_14773_ _14772_/X _26534_/Q _14773_/S vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19300_ _26829_/Q _26797_/Q _26765_/Q _26733_/Q _19297_/X _18930_/A vssd1 vssd1 vccd1
+ vccd1 _19300_/X sky130_fd_sc_hd__mux4_2
X_16512_ _16816_/A _16512_/B vssd1 vssd1 vccd1 vccd1 _16629_/B sky130_fd_sc_hd__xnor2_2
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13724_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17492_ _27429_/Q vssd1 vssd1 vccd1 vccd1 _17492_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19231_ _26954_/Q _26922_/Q _26890_/Q _26858_/Q _19208_/X _19116_/X vssd1 vssd1 vccd1
+ vccd1 _19231_/X sky130_fd_sc_hd__mux4_2
XFILLER_189_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16443_ _27388_/Q _16094_/A _16098_/A _25956_/Q _16442_/Y vssd1 vssd1 vccd1 vccd1
+ _16780_/B sky130_fd_sc_hd__a221o_1
X_13655_ _26913_/Q _13653_/X _13642_/X _13654_/Y vssd1 vssd1 vccd1 vccd1 _26913_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_182_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19162_ _27806_/Q _26567_/Q _26439_/Q _26119_/Q _19118_/X _19019_/X vssd1 vssd1 vccd1
+ vccd1 _19162_/X sky130_fd_sc_hd__mux4_2
X_13586_ _13602_/A vssd1 vssd1 vccd1 vccd1 _13670_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16374_ _16374_/A vssd1 vssd1 vccd1 vccd1 _16375_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18113_ _26148_/Q _26084_/Q _27012_/Q _26980_/Q _18041_/X _18112_/X vssd1 vssd1 vccd1
+ vccd1 _18114_/A sky130_fd_sc_hd__mux4_1
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15325_ _15325_/A vssd1 vssd1 vccd1 vccd1 _26302_/D sky130_fd_sc_hd__clkbuf_1
X_19093_ _19438_/A vssd1 vssd1 vccd1 vccd1 _19211_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18044_ _18358_/A vssd1 vssd1 vccd1 vccd1 _18044_/X sky130_fd_sc_hd__clkbuf_4
X_15256_ _14804_/X _26332_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15257_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14207_ _14220_/A vssd1 vssd1 vccd1 vccd1 _14207_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15187_ _15187_/A vssd1 vssd1 vccd1 vccd1 _26363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_513 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14138_ _14403_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14138_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19995_ _25641_/A vssd1 vssd1 vccd1 vccd1 _20340_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14069_ _26776_/Q _14058_/X _14064_/X _14068_/Y vssd1 vssd1 vccd1 vccd1 _26776_/D
+ sky130_fd_sc_hd__a31o_1
X_18946_ _19438_/A vssd1 vssd1 vccd1 vccd1 _19047_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18877_ _27795_/Q _26556_/Q _26428_/Q _26108_/Q _18793_/X _18851_/X vssd1 vssd1 vccd1
+ vccd1 _18877_/X sky130_fd_sc_hd__mux4_2
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17828_ _17828_/A _17827_/X vssd1 vssd1 vccd1 vccd1 _17828_/X sky130_fd_sc_hd__or2b_1
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ _17759_/A vssd1 vssd1 vccd1 vccd1 _25937_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20770_ _20770_/A vssd1 vssd1 vccd1 vccd1 _20770_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19429_ _26835_/Q _26803_/Q _26771_/Q _26739_/Q _19338_/X _19407_/X vssd1 vssd1 vccd1
+ vccd1 _19430_/B sky130_fd_sc_hd__mux4_1
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22440_ _22508_/A vssd1 vssd1 vccd1 vccd1 _22440_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22371_ _22457_/A vssd1 vssd1 vccd1 vccd1 _22436_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24110_ _24110_/A vssd1 vssd1 vccd1 vccd1 _27329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21322_ _21389_/A vssd1 vssd1 vccd1 vccd1 _21322_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25090_ _27976_/A _25089_/X _25104_/S vssd1 vssd1 vccd1 vccd1 _25091_/A sky130_fd_sc_hd__mux2_1
XFILLER_135_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24041_ _27096_/Q _23860_/A _23861_/A _27128_/Q _23862_/A vssd1 vssd1 vccd1 vccd1
+ _24041_/X sky130_fd_sc_hd__a221o_1
X_21253_ _21301_/A vssd1 vssd1 vccd1 vccd1 _21253_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_618 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20204_ _20236_/A vssd1 vssd1 vccd1 vccd1 _20204_/X sky130_fd_sc_hd__clkbuf_2
X_21184_ _21200_/A vssd1 vssd1 vccd1 vccd1 _21184_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27800_ _25650_/X _27800_/D vssd1 vssd1 vccd1 vccd1 _27800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20135_ _20151_/A vssd1 vssd1 vccd1 vccd1 _20135_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25992_ _26024_/CLK _25992_/D vssd1 vssd1 vccd1 vccd1 _25992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27731_ _27744_/CLK _27731_/D vssd1 vssd1 vccd1 vccd1 _27731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20066_ _20060_/X _20061_/X _20062_/X _20063_/X _20064_/X _20065_/X vssd1 vssd1 vccd1
+ vccd1 _20067_/A sky130_fd_sc_hd__mux4_1
X_24943_ _24947_/B _24943_/B vssd1 vssd1 vccd1 vccd1 _24944_/B sky130_fd_sc_hd__or2_1
XFILLER_100_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27662_ _27663_/CLK _27662_/D vssd1 vssd1 vccd1 vccd1 _27662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24874_ _24880_/C _24874_/B vssd1 vssd1 vccd1 vccd1 _24875_/B sky130_fd_sc_hd__or2_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater270 _27488_/CLK vssd1 vssd1 vccd1 vccd1 _27589_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26613_ _21456_/X _26613_/D vssd1 vssd1 vccd1 vccd1 _26613_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater281 _27523_/CLK vssd1 vssd1 vccd1 vccd1 _27592_/CLK sky130_fd_sc_hd__clkbuf_1
X_23825_ _27785_/Q vssd1 vssd1 vccd1 vccd1 _24014_/A sky130_fd_sc_hd__buf_2
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater292 _27468_/CLK vssd1 vssd1 vccd1 vccd1 _27461_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_304 _17898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 _18876_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27593_ _27593_/CLK _27593_/D vssd1 vssd1 vccd1 vccd1 _27593_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _24925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_337 _13204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 _16033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26544_ _21210_/X _26544_/D vssd1 vssd1 vccd1 vccd1 _26544_/Q sky130_fd_sc_hd__dfxtp_1
X_23756_ _27066_/Q _27098_/Q _23796_/S vssd1 vssd1 vccd1 vccd1 _23756_/X sky130_fd_sc_hd__mux2_1
X_20968_ _20968_/A vssd1 vssd1 vccd1 vccd1 _20968_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_359 _14791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22707_ _22697_/X _22698_/X _22699_/X _22700_/X _22702_/X _22704_/X vssd1 vssd1 vccd1
+ vccd1 _22708_/A sky130_fd_sc_hd__mux4_1
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23687_ _23687_/A vssd1 vssd1 vccd1 vccd1 _27248_/D sky130_fd_sc_hd__clkbuf_1
X_26475_ _20982_/X _26475_/D vssd1 vssd1 vccd1 vccd1 _26475_/Q sky130_fd_sc_hd__dfxtp_1
X_20899_ _20886_/X _20888_/X _20890_/X _20892_/X _20893_/X _20894_/X vssd1 vssd1 vccd1
+ vccd1 _20900_/A sky130_fd_sc_hd__mux4_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _27364_/Q _13108_/A _13082_/X _27332_/Q _13065_/X vssd1 vssd1 vccd1 vccd1
+ _14425_/A sky130_fd_sc_hd__a221oi_4
X_22638_ _22686_/A vssd1 vssd1 vccd1 vccd1 _22638_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25426_ _27751_/Q input64/X _25428_/S vssd1 vssd1 vccd1 vccd1 _25427_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28023__489 vssd1 vssd1 vccd1 vccd1 _28023__489/HI _28023_/A sky130_fd_sc_hd__conb_1
XFILLER_55_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25357_ _27720_/Q _25139_/A _25356_/Y _13423_/X vssd1 vssd1 vccd1 vccd1 _27720_/D
+ sky130_fd_sc_hd__o211a_1
X_13371_ _26986_/Q _13369_/X _13383_/S vssd1 vssd1 vccd1 vccd1 _13372_/A sky130_fd_sc_hd__mux2_1
X_22569_ _22561_/X _22562_/X _22563_/X _22564_/X _22565_/X _22566_/X vssd1 vssd1 vccd1
+ vccd1 _22570_/A sky130_fd_sc_hd__mux4_1
XFILLER_139_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15110_ _14801_/X _26397_/Q _15112_/S vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24308_ _24308_/A _24384_/B vssd1 vssd1 vccd1 vccd1 _27437_/D sky130_fd_sc_hd__nor2_1
X_16090_ _16639_/A _25907_/Q vssd1 vssd1 vccd1 vccd1 _16091_/A sky130_fd_sc_hd__or2_1
XFILLER_154_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25288_ _27508_/Q _27507_/Q _25347_/A vssd1 vssd1 vccd1 vccd1 _25288_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_957 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15041_ _15779_/A _15043_/B vssd1 vssd1 vccd1 vccd1 _15041_/Y sky130_fd_sc_hd__nor2_1
X_27027_ _22902_/X _27027_/D vssd1 vssd1 vccd1 vccd1 _27027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24239_ _24330_/A vssd1 vssd1 vccd1 vccd1 _24250_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_170_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18800_ _19448_/A vssd1 vssd1 vccd1 vccd1 _19324_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19780_ _19812_/A vssd1 vssd1 vccd1 vccd1 _19780_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16992_ _17338_/A vssd1 vssd1 vccd1 vccd1 _16992_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _26027_/Q _17731_/X _18735_/S vssd1 vssd1 vccd1 vccd1 _18732_/A sky130_fd_sc_hd__mux2_1
X_15943_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15943_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27929_ _27929_/A _15957_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18662_ _18662_/A vssd1 vssd1 vccd1 vccd1 _25996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15874_/Y sky130_fd_sc_hd__inv_2
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17613_ _17613_/A vssd1 vssd1 vccd1 vccd1 _25879_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _14825_/A vssd1 vssd1 vccd1 vccd1 _26517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _25437_/A vssd1 vssd1 vccd1 vccd1 _18594_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _17544_/A vssd1 vssd1 vccd1 vccd1 _25848_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ _14756_/A vssd1 vssd1 vccd1 vccd1 _14756_/X sky130_fd_sc_hd__buf_2
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _26895_/Q _13697_/X _13705_/X _13706_/Y vssd1 vssd1 vccd1 vccd1 _26895_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17475_ _17475_/A vssd1 vssd1 vccd1 vccd1 _25826_/D sky130_fd_sc_hd__clkbuf_1
X_14687_ _26563_/Q _14685_/X _14679_/X _14686_/Y vssd1 vssd1 vccd1 vccd1 _26563_/D
+ sky130_fd_sc_hd__a31o_1
X_19214_ _26537_/Q _26505_/Q _26473_/Q _27049_/Q _18926_/A _18923_/X vssd1 vssd1 vccd1
+ vccd1 _19214_/X sky130_fd_sc_hd__mux4_1
X_16426_ _16426_/A _16490_/B vssd1 vssd1 vccd1 vccd1 _16426_/Y sky130_fd_sc_hd__nor2_1
X_13638_ _26919_/Q _13626_/X _13629_/X _13637_/Y vssd1 vssd1 vccd1 vccd1 _26919_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19145_ _26278_/Q _26246_/Q _26214_/Q _26182_/Q _19144_/X _19074_/X vssd1 vssd1 vccd1
+ vccd1 _19145_/X sky130_fd_sc_hd__mux4_1
X_16357_ _16357_/A vssd1 vssd1 vccd1 vccd1 _16764_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13569_ _13934_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13569_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _15319_/A vssd1 vssd1 vccd1 vccd1 _15317_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19076_ _19488_/A vssd1 vssd1 vccd1 vccd1 _19076_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16288_ _27397_/Q _16297_/B vssd1 vssd1 vccd1 vccd1 _16288_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18027_ _18019_/X _18022_/X _18025_/X _18026_/X _17990_/X vssd1 vssd1 vccd1 vccd1
+ _18028_/C sky130_fd_sc_hd__a221o_1
X_15239_ _14779_/X _26340_/Q _15245_/S vssd1 vssd1 vccd1 vccd1 _15240_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19978_ _19972_/X _19973_/X _19974_/X _19975_/X _19976_/X _19977_/X vssd1 vssd1 vccd1
+ vccd1 _19979_/A sky130_fd_sc_hd__mux4_1
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18929_ _18929_/A vssd1 vssd1 vccd1 vccd1 _18929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21940_ _21940_/A vssd1 vssd1 vccd1 vccd1 _21940_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21871_ _21863_/X _21864_/X _21865_/X _21866_/X _21867_/X _21868_/X vssd1 vssd1 vccd1
+ vccd1 _21872_/A sky130_fd_sc_hd__mux4_1
XFILLER_131_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23610_ _23610_/A vssd1 vssd1 vccd1 vccd1 _27222_/D sky130_fd_sc_hd__clkbuf_1
X_20822_ _20816_/X _20817_/X _20818_/X _20819_/X _20820_/X _20821_/X vssd1 vssd1 vccd1
+ vccd1 _20823_/A sky130_fd_sc_hd__mux4_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24590_ _27655_/Q _24598_/B vssd1 vssd1 vccd1 vccd1 _24591_/A sky130_fd_sc_hd__and2_1
XFILLER_36_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23541_ _23541_/A vssd1 vssd1 vccd1 vccd1 _27203_/D sky130_fd_sc_hd__clkbuf_1
X_20753_ _20753_/A vssd1 vssd1 vccd1 vccd1 _20753_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26260_ _20223_/X _26260_/D vssd1 vssd1 vccd1 vccd1 _26260_/Q sky130_fd_sc_hd__dfxtp_1
X_23472_ _23485_/A vssd1 vssd1 vccd1 vccd1 _23483_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_196_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20684_ _20684_/A vssd1 vssd1 vccd1 vccd1 _20684_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25211_ _25211_/A _25211_/B vssd1 vssd1 vccd1 vccd1 _25212_/B sky130_fd_sc_hd__nand2_1
X_22423_ _22417_/X _22418_/X _22419_/X _22420_/X _22421_/X _22422_/X vssd1 vssd1 vccd1
+ vccd1 _22424_/A sky130_fd_sc_hd__mux4_1
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26191_ _19981_/X _26191_/D vssd1 vssd1 vccd1 vccd1 _26191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25142_ _25308_/A vssd1 vssd1 vccd1 vccd1 _25142_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22354_ _22422_/A vssd1 vssd1 vccd1 vccd1 _22354_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21305_ _22613_/A vssd1 vssd1 vccd1 vccd1 _21651_/A sky130_fd_sc_hd__clkbuf_2
X_25073_ _27077_/Q _27109_/Q _25088_/S vssd1 vssd1 vccd1 vccd1 _25073_/X sky130_fd_sc_hd__mux2_1
X_22285_ _22457_/A vssd1 vssd1 vccd1 vccd1 _22350_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24024_ _24022_/X _24023_/X _24031_/S vssd1 vssd1 vccd1 vccd1 _24024_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21236_ _21583_/A vssd1 vssd1 vccd1 vccd1 _21303_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21167_ _21199_/A vssd1 vssd1 vccd1 vccd1 _21167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20118_ _20150_/A vssd1 vssd1 vccd1 vccd1 _20118_/X sky130_fd_sc_hd__clkbuf_2
X_21098_ _21114_/A vssd1 vssd1 vccd1 vccd1 _21098_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25975_ _26056_/CLK _25975_/D vssd1 vssd1 vccd1 vccd1 _25975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27714_ _27716_/CLK _27714_/D vssd1 vssd1 vccd1 vccd1 _27714_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _27824_/Q _25297_/A vssd1 vssd1 vccd1 vccd1 _12941_/A sky130_fd_sc_hd__and2_1
X_20049_ _20065_/A vssd1 vssd1 vccd1 vccd1 _20049_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24926_ _24925_/B _24925_/C _24925_/A vssd1 vssd1 vccd1 vccd1 _24927_/B sky130_fd_sc_hd__a21oi_1
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27645_ _27645_/CLK _27645_/D vssd1 vssd1 vccd1 vccd1 _27645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24857_ _27761_/Q _24857_/B vssd1 vssd1 vccd1 vccd1 _24858_/B sky130_fd_sc_hd__nor2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _19336_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _20589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_123 _22546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _15771_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14610_/Y sky130_fd_sc_hd__nor2_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _25066_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23808_ _24046_/S vssd1 vssd1 vccd1 vccd1 _23845_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15590_ _15590_/A vssd1 vssd1 vccd1 vccd1 _26185_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27576_ _27576_/CLK _27576_/D vssd1 vssd1 vccd1 vccd1 _27576_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24788_ _27628_/Q _24785_/X _24786_/Y _24787_/X vssd1 vssd1 vccd1 vccd1 _27628_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _13056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _13347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_167 _13408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_178 _16289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14541_ _26616_/Q _14530_/X _14536_/X _14540_/Y vssd1 vssd1 vccd1 vccd1 _26616_/D
+ sky130_fd_sc_hd__a31o_1
X_26527_ _21158_/X _26527_/D vssd1 vssd1 vccd1 vccd1 _26527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _16495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23739_ _23990_/A vssd1 vssd1 vccd1 vccd1 _23849_/A sky130_fd_sc_hd__buf_2
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17260_ _17258_/X _17259_/X _17296_/S vssd1 vssd1 vccd1 vccd1 _17260_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14472_ _15738_/A _14483_/B vssd1 vssd1 vccd1 vccd1 _14472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26458_ _20918_/X _26458_/D vssd1 vssd1 vccd1 vccd1 _26458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16211_ _17420_/B _16233_/B vssd1 vssd1 vccd1 vccd1 _16211_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13423_ _25733_/B vssd1 vssd1 vccd1 vccd1 _13423_/X sky130_fd_sc_hd__buf_4
X_25409_ _27743_/Q input55/X _25413_/S vssd1 vssd1 vccd1 vccd1 _25410_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17191_ _17252_/A vssd1 vssd1 vccd1 vccd1 _17191_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26389_ _20667_/X _26389_/D vssd1 vssd1 vccd1 vccd1 _26389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16142_ _16796_/A vssd1 vssd1 vccd1 vccd1 _16833_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ _13421_/S vssd1 vssd1 vccd1 vccd1 _13367_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16073_ _16623_/A _16845_/B _16073_/C vssd1 vssd1 vccd1 vccd1 _16602_/A sky130_fd_sc_hd__and3_1
XFILLER_6_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13285_ _27017_/Q _13150_/X _13291_/S vssd1 vssd1 vccd1 vccd1 _13286_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15024_ _15762_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19901_ _19901_/A vssd1 vssd1 vccd1 vccd1 _19901_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19832_ _19832_/A vssd1 vssd1 vccd1 vccd1 _19899_/A sky130_fd_sc_hd__buf_2
XFILLER_2_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19763_ _19763_/A vssd1 vssd1 vccd1 vccd1 _19763_/X sky130_fd_sc_hd__clkbuf_1
X_16975_ _27608_/Q _24635_/A _16974_/Y _24522_/A _24633_/A vssd1 vssd1 vccd1 vccd1
+ _16976_/B sky130_fd_sc_hd__a32o_1
XFILLER_77_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18714_ _18714_/A vssd1 vssd1 vccd1 vccd1 _26019_/D sky130_fd_sc_hd__clkbuf_1
X_15926_ _15930_/A vssd1 vssd1 vccd1 vccd1 _15926_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19694_ _19726_/A vssd1 vssd1 vccd1 vccd1 _19694_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 io_in[8] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18645_ _18645_/A vssd1 vssd1 vccd1 vccd1 _25988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15857_ _15988_/A vssd1 vssd1 vccd1 vccd1 _15862_/A sky130_fd_sc_hd__buf_8
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _14807_/X _26523_/Q _14811_/S vssd1 vssd1 vccd1 vccd1 _14809_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18576_ _26297_/Q _26265_/Q _26233_/Q _26201_/Q _18004_/X _18481_/X vssd1 vssd1 vccd1
+ vccd1 _18576_/X sky130_fd_sc_hd__mux4_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15788_ _13058_/X _26104_/Q _15794_/S vssd1 vssd1 vccd1 vccd1 _15789_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17527_ _27378_/Q vssd1 vssd1 vccd1 vccd1 _25735_/B sky130_fd_sc_hd__clkbuf_2
X_14739_ _14739_/A vssd1 vssd1 vccd1 vccd1 _26545_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ _17456_/X _25821_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17459_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16409_ _16359_/A _16447_/C _16733_/B _16369_/X vssd1 vssd1 vccd1 vccd1 _16410_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_177_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ input9/X vssd1 vssd1 vccd1 vccd1 _20788_/A sky130_fd_sc_hd__inv_2
XFILLER_118_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19128_ _19126_/X _19127_/X _19173_/S vssd1 vssd1 vccd1 vccd1 _19128_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19059_ _19107_/A _19059_/B _19059_/C vssd1 vssd1 vccd1 vccd1 _19060_/A sky130_fd_sc_hd__and3_1
XFILLER_145_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22070_ _22086_/A vssd1 vssd1 vccd1 vccd1 _22070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1089 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21021_ _21007_/X _21008_/X _21009_/X _21010_/X _21011_/X _21012_/X vssd1 vssd1 vccd1
+ vccd1 _21022_/A sky130_fd_sc_hd__mux4_1
XFILLER_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25760_ _17456_/X _27836_/Q _25768_/S vssd1 vssd1 vccd1 vccd1 _25761_/A sky130_fd_sc_hd__mux2_1
X_22972_ _22972_/A vssd1 vssd1 vccd1 vccd1 _22972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24711_ _27186_/Q _24711_/B vssd1 vssd1 vccd1 vccd1 _24711_/X sky130_fd_sc_hd__or2_1
X_21923_ _21911_/X _21912_/X _21913_/X _21914_/X _21916_/X _21918_/X vssd1 vssd1 vccd1
+ vccd1 _21924_/A sky130_fd_sc_hd__mux4_1
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25691_ _25723_/A vssd1 vssd1 vccd1 vccd1 _25691_/X sky130_fd_sc_hd__clkbuf_1
X_27430_ _27430_/CLK _27430_/D vssd1 vssd1 vccd1 vccd1 _27430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21854_ _21854_/A vssd1 vssd1 vccd1 vccd1 _21854_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24642_ _24841_/A vssd1 vssd1 vccd1 vccd1 _24700_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20805_ _20853_/A vssd1 vssd1 vccd1 vccd1 _20805_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27361_ _27473_/CLK _27361_/D vssd1 vssd1 vccd1 vccd1 _27361_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21785_ _21777_/X _21778_/X _21779_/X _21780_/X _21781_/X _21782_/X vssd1 vssd1 vccd1
+ vccd1 _21786_/A sky130_fd_sc_hd__mux4_1
X_24573_ _24573_/A vssd1 vssd1 vccd1 vccd1 _27547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26312_ _20403_/X _26312_/D vssd1 vssd1 vccd1 vccd1 _26312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20736_ _20722_/X _20723_/X _20724_/X _20725_/X _20726_/X _20727_/X vssd1 vssd1 vccd1
+ vccd1 _20737_/A sky130_fd_sc_hd__mux4_1
X_23524_ _27757_/Q vssd1 vssd1 vccd1 vccd1 _24835_/A sky130_fd_sc_hd__buf_2
X_27292_ _27293_/CLK _27292_/D vssd1 vssd1 vccd1 vccd1 _27292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26243_ _20159_/X _26243_/D vssd1 vssd1 vccd1 vccd1 _26243_/Q sky130_fd_sc_hd__dfxtp_1
X_23455_ _23482_/A vssd1 vssd1 vccd1 vccd1 _23455_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20667_ _20667_/A vssd1 vssd1 vccd1 vccd1 _20667_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22406_ _22422_/A vssd1 vssd1 vccd1 vccd1 _22406_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23386_ _24862_/A _23383_/Y _27256_/Q _24794_/A _23385_/X vssd1 vssd1 vccd1 vccd1
+ _23393_/B sky130_fd_sc_hd__a221o_1
XFILLER_52_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26174_ _19915_/X _26174_/D vssd1 vssd1 vccd1 vccd1 _26174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20598_ _20598_/A vssd1 vssd1 vccd1 vccd1 _20598_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_457 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22337_ _22331_/X _22332_/X _22333_/X _22334_/X _22335_/X _22336_/X vssd1 vssd1 vccd1
+ vccd1 _22338_/A sky130_fd_sc_hd__mux4_1
X_25125_ _27522_/Q _27490_/Q vssd1 vssd1 vccd1 vccd1 _25127_/A sky130_fd_sc_hd__and2_1
XFILLER_87_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25056_ _25102_/S vssd1 vssd1 vccd1 vccd1 _25088_/S sky130_fd_sc_hd__clkbuf_2
X_13070_ _27299_/Q _13169_/B vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__and2_1
X_22268_ _22336_/A vssd1 vssd1 vccd1 vccd1 _22268_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24007_ _27852_/Q _27156_/Q _25901_/Q _25869_/Q _23967_/X _23991_/X vssd1 vssd1 vccd1
+ vccd1 _24007_/X sky130_fd_sc_hd__mux4_1
X_21219_ _21211_/X _21212_/X _21213_/X _21214_/X _21216_/X _21218_/X vssd1 vssd1 vccd1
+ vccd1 _21220_/A sky130_fd_sc_hd__mux4_1
XFILLER_2_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22199_ _22457_/A vssd1 vssd1 vccd1 vccd1 _22264_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16760_ _25945_/Q _16375_/B _16563_/B _14527_/A vssd1 vssd1 vccd1 vccd1 _16761_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_98_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ _26803_/Q _13969_/X _13965_/X _13971_/Y vssd1 vssd1 vccd1 vccd1 _26803_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25958_ _25958_/CLK _25958_/D vssd1 vssd1 vccd1 vccd1 _25958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15711_ _26133_/Q _15705_/X _15697_/X _15710_/Y vssd1 vssd1 vccd1 vccd1 _26133_/D
+ sky130_fd_sc_hd__a31o_1
X_12923_ input61/X input62/X input64/X input65/X vssd1 vssd1 vccd1 vccd1 _12929_/C
+ sky130_fd_sc_hd__nand4_1
X_24909_ _24935_/A vssd1 vssd1 vccd1 vccd1 _24909_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16691_ _16686_/Y _16687_/X _16690_/X vssd1 vssd1 vccd1 vccd1 _24235_/A sky130_fd_sc_hd__a21oi_1
X_25889_ _27144_/CLK _25889_/D vssd1 vssd1 vccd1 vccd1 _25889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18430_ _26834_/Q _26802_/Q _26770_/Q _26738_/Q _18358_/X _18380_/X vssd1 vssd1 vccd1
+ vccd1 _18430_/X sky130_fd_sc_hd__mux4_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27628_ _27629_/CLK _27628_/D vssd1 vssd1 vccd1 vccd1 _27628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15642_ _15642_/A vssd1 vssd1 vccd1 vccd1 _26162_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _26703_/Q _26671_/Q _26639_/Q _26607_/Q _18360_/X _18249_/X vssd1 vssd1 vccd1
+ vccd1 _18362_/A sky130_fd_sc_hd__mux4_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27559_ _27559_/CLK _27559_/D vssd1 vssd1 vccd1 vccd1 _27559_/Q sky130_fd_sc_hd__dfxtp_1
X_15573_ _26192_/Q _14740_/A _15573_/S vssd1 vssd1 vccd1 vccd1 _15574_/A sky130_fd_sc_hd__mux2_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _17312_/A vssd1 vssd1 vccd1 vccd1 _27940_/A sky130_fd_sc_hd__clkbuf_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14524_ _14524_/A vssd1 vssd1 vccd1 vccd1 _15777_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18292_ _26700_/Q _26668_/Q _26636_/Q _26604_/Q _18004_/X _18005_/X vssd1 vssd1 vccd1
+ vccd1 _18293_/A sky130_fd_sc_hd__mux4_2
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17243_ _25830_/Q _26029_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17243_/X sky130_fd_sc_hd__mux2_1
X_14455_ _14510_/A vssd1 vssd1 vccd1 vccd1 _14455_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ _26975_/Q _13405_/X _13415_/S vssd1 vssd1 vccd1 vccd1 _13407_/A sky130_fd_sc_hd__mux2_1
X_17174_ _17172_/X _17173_/X _17174_/S vssd1 vssd1 vccd1 vccd1 _17174_/X sky130_fd_sc_hd__mux2_2
X_14386_ _14386_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _14386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ _16845_/A _16125_/B vssd1 vssd1 vccd1 vccd1 _16304_/A sky130_fd_sc_hd__and2_1
X_13337_ _14727_/A vssd1 vssd1 vccd1 vccd1 _13337_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16056_ _27475_/Q vssd1 vssd1 vccd1 vccd1 _16056_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13268_ _13268_/A vssd1 vssd1 vccd1 vccd1 _27025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15007_ _26441_/Q _15002_/X _15003_/X _15006_/Y vssd1 vssd1 vccd1 vccd1 _26441_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _27041_/Q _13198_/X _13199_/S vssd1 vssd1 vccd1 vccd1 _13200_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19815_ _19815_/A vssd1 vssd1 vccd1 vccd1 _19815_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16958_ _27584_/Q _24626_/D vssd1 vssd1 vccd1 vccd1 _24636_/B sky130_fd_sc_hd__nor2_1
XFILLER_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19746_ _19832_/A vssd1 vssd1 vccd1 vccd1 _19813_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15909_ _15912_/A vssd1 vssd1 vccd1 vccd1 _15909_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19677_ _19677_/A vssd1 vssd1 vccd1 vccd1 _19677_/X sky130_fd_sc_hd__clkbuf_1
X_16889_ _16887_/X _16797_/X _16888_/Y _16877_/X vssd1 vssd1 vccd1 vccd1 _24256_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18628_ _25981_/Q _17686_/X _18630_/S vssd1 vssd1 vccd1 vccd1 _18629_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18559_ _17886_/S _18558_/X _18483_/X vssd1 vssd1 vccd1 vccd1 _18559_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21570_ _21570_/A vssd1 vssd1 vccd1 vccd1 _21570_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_12 _25888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _27141_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ _20521_/A vssd1 vssd1 vccd1 vccd1 _20521_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_34 _17723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_45 _17923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 _18221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23240_ _17504_/X _27155_/Q _23248_/S vssd1 vssd1 vccd1 vccd1 _23241_/A sky130_fd_sc_hd__mux2_1
XANTENNA_67 _18339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20452_ _20500_/A vssd1 vssd1 vccd1 vccd1 _20452_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_78 _18557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 _18943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23171_ _23171_/A vssd1 vssd1 vccd1 vccd1 _27124_/D sky130_fd_sc_hd__clkbuf_1
X_20383_ _20383_/A vssd1 vssd1 vccd1 vccd1 _20383_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22122_ _22122_/A vssd1 vssd1 vccd1 vccd1 _22122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22053_ _22085_/A vssd1 vssd1 vccd1 vccd1 _22053_/X sky130_fd_sc_hd__clkbuf_1
X_26930_ _22568_/X _26930_/D vssd1 vssd1 vccd1 vccd1 _26930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21004_ _21004_/A vssd1 vssd1 vccd1 vccd1 _21004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26861_ _22324_/X _26861_/D vssd1 vssd1 vccd1 vccd1 _26861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25812_ _26012_/CLK _25812_/D vssd1 vssd1 vccd1 vccd1 _25812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26792_ _22078_/X _26792_/D vssd1 vssd1 vccd1 vccd1 _26792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25743_ _25743_/A vssd1 vssd1 vccd1 vccd1 _27828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22955_ _22955_/A vssd1 vssd1 vccd1 vccd1 _22955_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21906_ _21906_/A vssd1 vssd1 vccd1 vccd1 _21906_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25674_ _25722_/A vssd1 vssd1 vccd1 vccd1 _25674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22886_ _22886_/A vssd1 vssd1 vccd1 vccd1 _22886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27413_ _27413_/CLK _27413_/D vssd1 vssd1 vccd1 vccd1 _27413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24625_ _24625_/A vssd1 vssd1 vccd1 vccd1 _27571_/D sky130_fd_sc_hd__clkbuf_1
X_21837_ _21825_/X _21826_/X _21827_/X _21828_/X _21830_/X _21832_/X vssd1 vssd1 vccd1
+ vccd1 _21838_/A sky130_fd_sc_hd__mux4_1
XFILLER_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27344_ _27559_/CLK _27344_/D vssd1 vssd1 vccd1 vccd1 _27344_/Q sky130_fd_sc_hd__dfxtp_2
X_21768_ _21768_/A vssd1 vssd1 vccd1 vccd1 _21768_/X sky130_fd_sc_hd__clkbuf_1
X_24556_ _24589_/A vssd1 vssd1 vccd1 vccd1 _24565_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_491 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20719_ _20719_/A vssd1 vssd1 vccd1 vccd1 _20719_/X sky130_fd_sc_hd__clkbuf_1
X_23507_ _23507_/A _23507_/B vssd1 vssd1 vccd1 vccd1 _23600_/A sky130_fd_sc_hd__or2_4
XFILLER_54_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27275_ _27278_/CLK _27275_/D vssd1 vssd1 vccd1 vccd1 _27275_/Q sky130_fd_sc_hd__dfxtp_1
X_21699_ _21689_/X _21690_/X _21691_/X _21692_/X _21693_/X _21694_/X vssd1 vssd1 vccd1
+ vccd1 _21700_/A sky130_fd_sc_hd__mux4_1
XFILLER_169_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24487_ _24636_/A vssd1 vssd1 vccd1 vccd1 _24631_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ _15335_/A _14534_/B vssd1 vssd1 vccd1 vccd1 _14257_/A sky130_fd_sc_hd__nand2b_1
X_26226_ _20107_/X _26226_/D vssd1 vssd1 vccd1 vccd1 _26226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23438_ _27169_/Q _23443_/B vssd1 vssd1 vccd1 vccd1 _23438_/X sky130_fd_sc_hd__or2_1
XFILLER_109_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14171_ _26739_/Q _14157_/X _14167_/X _14170_/Y vssd1 vssd1 vccd1 vccd1 _26739_/D
+ sky130_fd_sc_hd__a31o_1
X_23369_ _27766_/Q vssd1 vssd1 vccd1 vccd1 _24767_/A sky130_fd_sc_hd__inv_2
X_26157_ _19861_/X _26157_/D vssd1 vssd1 vccd1 vccd1 _26157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25108_ _25108_/A _25733_/A vssd1 vssd1 vccd1 vccd1 _25108_/Y sky130_fd_sc_hd__nand2_1
X_13122_ _14747_/A vssd1 vssd1 vccd1 vccd1 _13122_/X sky130_fd_sc_hd__buf_2
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26088_ _19618_/X _26088_/D vssd1 vssd1 vccd1 vccd1 _26088_/Q sky130_fd_sc_hd__dfxtp_1
X_17930_ _17930_/A _17813_/X vssd1 vssd1 vccd1 vccd1 _17930_/X sky130_fd_sc_hd__or2b_1
XFILLER_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13053_ _13053_/A vssd1 vssd1 vccd1 vccd1 _27065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25039_ _27073_/Q _27105_/Q _25047_/S vssd1 vssd1 vccd1 vccd1 _25039_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17861_ _26939_/Q _26907_/Q _26875_/Q _26843_/Q _17789_/X _17791_/X vssd1 vssd1 vccd1
+ vccd1 _17861_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16812_ _16812_/A _16812_/B vssd1 vssd1 vccd1 vccd1 _16844_/A sky130_fd_sc_hd__nand2_1
X_19600_ _19600_/A vssd1 vssd1 vccd1 vccd1 _19600_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17792_ _26938_/Q _26906_/Q _26874_/Q _26842_/Q _17789_/X _17791_/X vssd1 vssd1 vccd1
+ vccd1 _17792_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19531_ _19567_/A _19531_/B _19531_/C vssd1 vssd1 vccd1 vccd1 _19532_/A sky130_fd_sc_hd__and3_1
X_16743_ _16747_/A _16743_/B vssd1 vssd1 vccd1 vccd1 _16743_/Y sky130_fd_sc_hd__nand2_1
X_13955_ _26807_/Q _13949_/X _13944_/X _13954_/Y vssd1 vssd1 vccd1 vccd1 _26807_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19462_ _19524_/A _19462_/B vssd1 vssd1 vccd1 vccd1 _19462_/X sky130_fd_sc_hd__or2_1
X_16674_ _16674_/A vssd1 vssd1 vccd1 vccd1 _16852_/A sky130_fd_sc_hd__clkbuf_1
X_13886_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18413_ _18311_/X _18406_/X _18411_/X _18412_/X vssd1 vssd1 vccd1 vccd1 _18423_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _15693_/S vssd1 vssd1 vccd1 vccd1 _15634_/S sky130_fd_sc_hd__clkbuf_2
X_19393_ _19393_/A vssd1 vssd1 vccd1 vccd1 _19393_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _18344_/A _18020_/A vssd1 vssd1 vccd1 vccd1 _18344_/X sky130_fd_sc_hd__or2b_1
XFILLER_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _26200_/Q _14715_/A _15562_/S vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14507_/A vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__clkbuf_2
X_18275_ _18198_/X _18272_/X _18274_/X _18203_/X vssd1 vssd1 vccd1 vccd1 _18275_/X
+ sky130_fd_sc_hd__o211a_1
X_15487_ _15487_/A vssd1 vssd1 vccd1 vccd1 _26231_/D sky130_fd_sc_hd__clkbuf_1
X_17226_ _17226_/A vssd1 vssd1 vccd1 vccd1 _27933_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_175_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14438_ _14438_/A vssd1 vssd1 vccd1 vccd1 _15714_/A sky130_fd_sc_hd__buf_2
Xinput10 la1_data_in[10] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
Xinput21 la1_data_in[20] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 la1_data_in[30] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_2
Xinput43 la1_oenb[11] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_6
Xinput54 la1_oenb[21] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_4
X_17157_ _17155_/X _17157_/B vssd1 vssd1 vccd1 vccd1 _17157_/X sky130_fd_sc_hd__and2b_1
X_14369_ _14369_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14369_/Y sky130_fd_sc_hd__nor2_1
Xinput65 la1_oenb[31] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_4
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16108_ _16108_/A vssd1 vssd1 vccd1 vccd1 _16109_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17088_ _17052_/X _17082_/X _17085_/X _17087_/X vssd1 vssd1 vccd1 vccd1 _17088_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16039_ _27476_/Q _27475_/Q _27474_/Q vssd1 vssd1 vccd1 vccd1 _16062_/B sky130_fd_sc_hd__or3_1
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19729_ _19729_/A vssd1 vssd1 vccd1 vccd1 _19729_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22740_ _22772_/A vssd1 vssd1 vccd1 vccd1 _22740_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22671_ _22665_/X _22666_/X _22667_/X _22668_/X _22669_/X _22670_/X vssd1 vssd1 vccd1
+ vccd1 _22672_/A sky130_fd_sc_hd__mux4_1
XFILLER_164_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21622_ _21622_/A vssd1 vssd1 vccd1 vccd1 _21622_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24410_ _24410_/A vssd1 vssd1 vccd1 vccd1 _27484_/D sky130_fd_sc_hd__clkbuf_1
X_25390_ _25390_/A vssd1 vssd1 vccd1 vccd1 _27734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21553_ _21545_/X _21546_/X _21547_/X _21548_/X _21549_/X _21550_/X vssd1 vssd1 vccd1
+ vccd1 _21554_/A sky130_fd_sc_hd__mux4_1
X_24341_ _24363_/A vssd1 vssd1 vccd1 vccd1 _24350_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_194_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20504_ _20496_/X _20497_/X _20498_/X _20499_/X _20500_/X _20501_/X vssd1 vssd1 vccd1
+ vccd1 _20505_/A sky130_fd_sc_hd__mux4_1
XFILLER_53_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24272_ _16188_/X _16190_/Y _16191_/X _24269_/X vssd1 vssd1 vccd1 vccd1 _27410_/D
+ sky130_fd_sc_hd__o31a_1
X_27060_ _23016_/X _27060_/D vssd1 vssd1 vccd1 vccd1 _27060_/Q sky130_fd_sc_hd__dfxtp_1
X_21484_ _21484_/A vssd1 vssd1 vccd1 vccd1 _21484_/X sky130_fd_sc_hd__clkbuf_1
X_23223_ _23223_/A vssd1 vssd1 vccd1 vccd1 _27147_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26011_ _27676_/CLK _26011_/D vssd1 vssd1 vccd1 vccd1 _26011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20435_ _20435_/A vssd1 vssd1 vccd1 vccd1 _20435_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23154_ _27117_/Q _17737_/X _23154_/S vssd1 vssd1 vccd1 vccd1 _23155_/A sky130_fd_sc_hd__mux2_1
X_20366_ _20354_/X _20357_/X _20360_/X _20363_/X _20364_/X _20365_/X vssd1 vssd1 vccd1
+ vccd1 _20367_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22105_ _22453_/A vssd1 vssd1 vccd1 vccd1 _22174_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23085_ _23085_/A vssd1 vssd1 vccd1 vccd1 _27086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27962_ _27962_/A _15873_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_20297_ _20297_/A vssd1 vssd1 vccd1 vccd1 _20297_/X sky130_fd_sc_hd__clkbuf_1
X_22036_ _22084_/A vssd1 vssd1 vccd1 vccd1 _22036_/X sky130_fd_sc_hd__clkbuf_1
X_26913_ _22500_/X _26913_/D vssd1 vssd1 vccd1 vccd1 _26913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26844_ _22260_/X _26844_/D vssd1 vssd1 vccd1 vccd1 _26844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26775_ _22026_/X _26775_/D vssd1 vssd1 vccd1 vccd1 _26775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23987_ _23985_/X _23986_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23987_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ _13740_/A vssd1 vssd1 vccd1 vccd1 _13751_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25726_ _25726_/A vssd1 vssd1 vccd1 vccd1 _25726_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22938_ _22938_/A vssd1 vssd1 vccd1 vccd1 _22938_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _26906_/Q _13665_/X _13593_/B _13670_/Y vssd1 vssd1 vccd1 vccd1 _26906_/D
+ sky130_fd_sc_hd__a31o_1
X_25657_ _25657_/A vssd1 vssd1 vccd1 vccd1 _25723_/A sky130_fd_sc_hd__clkbuf_2
X_22869_ _22869_/A vssd1 vssd1 vccd1 vccd1 _22869_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15410_ _26265_/Q _13319_/X _15418_/S vssd1 vssd1 vccd1 vccd1 _15411_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24608_ _24608_/A vssd1 vssd1 vccd1 vccd1 _27563_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16390_ _16747_/A _16390_/B vssd1 vssd1 vccd1 vccd1 _16393_/B sky130_fd_sc_hd__xnor2_1
X_25588_ _24800_/A _25564_/X _25586_/X _25587_/Y _25557_/X vssd1 vssd1 vccd1 vccd1
+ _27778_/D sky130_fd_sc_hd__a221oi_1
XFILLER_197_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27327_ _27327_/CLK _27327_/D vssd1 vssd1 vccd1 vccd1 _27327_/Q sky130_fd_sc_hd__dfxtp_1
X_15341_ _15341_/A vssd1 vssd1 vccd1 vccd1 _26296_/D sky130_fd_sc_hd__clkbuf_1
X_24539_ _24534_/X _24386_/A _24545_/S vssd1 vssd1 vccd1 vccd1 _24540_/B sky130_fd_sc_hd__mux2_1
XFILLER_145_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18060_ _26690_/Q _26658_/Q _26626_/Q _26594_/Q _18036_/X _17928_/X vssd1 vssd1 vccd1
+ vccd1 _18061_/A sky130_fd_sc_hd__mux4_1
XFILLER_157_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27258_ _27258_/CLK _27258_/D vssd1 vssd1 vccd1 vccd1 _27258_/Q sky130_fd_sc_hd__dfxtp_1
X_15272_ _15272_/A vssd1 vssd1 vccd1 vccd1 _26326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17011_ _17387_/S vssd1 vssd1 vccd1 vccd1 _17067_/S sky130_fd_sc_hd__clkbuf_2
X_14223_ _14401_/A _14226_/B vssd1 vssd1 vccd1 vccd1 _14223_/Y sky130_fd_sc_hd__nor2_1
X_26209_ _20043_/X _26209_/D vssd1 vssd1 vccd1 vccd1 _26209_/Q sky130_fd_sc_hd__dfxtp_1
X_27189_ _27751_/CLK _27189_/D vssd1 vssd1 vccd1 vccd1 _27189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14154_ _26745_/Q _14142_/X _14151_/X _14153_/Y vssd1 vssd1 vccd1 vccd1 _26745_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ _14737_/A vssd1 vssd1 vccd1 vccd1 _13105_/X sky130_fd_sc_hd__buf_2
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14085_ _14350_/A _14085_/B vssd1 vssd1 vccd1 vccd1 _14085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18962_ _19391_/A vssd1 vssd1 vccd1 vccd1 _19057_/S sky130_fd_sc_hd__clkbuf_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17913_ _18012_/A vssd1 vssd1 vccd1 vccd1 _17913_/X sky130_fd_sc_hd__buf_4
X_13036_ _27302_/Q _13125_/B vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__and2_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18893_ _18893_/A vssd1 vssd1 vccd1 vccd1 _26044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17844_ _26522_/Q _26490_/Q _26458_/Q _27034_/Q _17841_/X _17843_/X vssd1 vssd1 vccd1
+ vccd1 _17844_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17775_ _27439_/Q vssd1 vssd1 vccd1 vccd1 _17775_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14987_ _26448_/Q _14974_/X _14976_/X _14986_/Y vssd1 vssd1 vccd1 vccd1 _26448_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19514_ _19514_/A vssd1 vssd1 vccd1 vccd1 _26070_/D sky130_fd_sc_hd__clkbuf_1
X_16726_ _16481_/A _16606_/Y _16450_/Y vssd1 vssd1 vccd1 vccd1 _16726_/Y sky130_fd_sc_hd__a21oi_1
X_13938_ _13938_/A _13940_/B vssd1 vssd1 vccd1 vccd1 _13938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19445_ _19445_/A vssd1 vssd1 vccd1 vccd1 _19445_/X sky130_fd_sc_hd__clkbuf_2
X_16657_ _16824_/A vssd1 vssd1 vccd1 vccd1 _16658_/A sky130_fd_sc_hd__inv_2
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13869_ _26838_/Q _13865_/X _13855_/X _13868_/Y vssd1 vssd1 vccd1 vccd1 _26838_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15608_ _15608_/A vssd1 vssd1 vccd1 vccd1 _15617_/S sky130_fd_sc_hd__clkbuf_2
X_19376_ _26160_/Q _26096_/Q _27024_/Q _26992_/Q _18807_/X _18810_/X vssd1 vssd1 vccd1
+ vccd1 _19377_/B sky130_fd_sc_hd__mux4_1
X_16588_ _16831_/B _16588_/B vssd1 vssd1 vccd1 vccd1 _16636_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18327_ _18279_/X _18325_/X _18326_/X vssd1 vssd1 vccd1 vccd1 _18327_/X sky130_fd_sc_hd__o21a_1
XFILLER_72_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _13210_/X _26207_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15540_/A sky130_fd_sc_hd__mux2_1
XFILLER_175_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _18162_/X _18257_/X _18211_/X vssd1 vssd1 vccd1 vccd1 _18258_/X sky130_fd_sc_hd__o21a_1
XFILLER_176_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _17181_/X _17208_/X _17159_/X vssd1 vssd1 vccd1 vccd1 _17209_/X sky130_fd_sc_hd__a21bo_1
XFILLER_191_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18189_ _18305_/A vssd1 vssd1 vccd1 vccd1 _18189_/X sky130_fd_sc_hd__buf_2
XFILLER_190_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20220_ _20236_/A vssd1 vssd1 vccd1 vccd1 _20220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20151_ _20151_/A vssd1 vssd1 vccd1 vccd1 _20151_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20082_ _20340_/A vssd1 vssd1 vccd1 vccd1 _20151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23910_ _27081_/Q _23907_/X _23908_/X _27113_/Q _23909_/X vssd1 vssd1 vccd1 vccd1
+ _23910_/X sky130_fd_sc_hd__a221o_1
XFILLER_112_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24890_ _24914_/A vssd1 vssd1 vccd1 vccd1 _24890_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater430 _25969_/CLK vssd1 vssd1 vccd1 vccd1 _26059_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23841_ _23800_/X _23839_/X _23840_/X _23816_/X vssd1 vssd1 vccd1 vccd1 _27279_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26560_ _21276_/X _26560_/D vssd1 vssd1 vccd1 vccd1 _26560_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _20984_/A vssd1 vssd1 vccd1 vccd1 _20984_/X sky130_fd_sc_hd__clkbuf_1
X_23772_ _23770_/X _23771_/X _23795_/S vssd1 vssd1 vccd1 vccd1 _23772_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25511_ _27702_/Q _25509_/X _25510_/X vssd1 vssd1 vccd1 vccd1 _25511_/Y sky130_fd_sc_hd__a21oi_1
X_22723_ _22771_/A vssd1 vssd1 vccd1 vccd1 _22723_/X sky130_fd_sc_hd__clkbuf_2
X_26491_ _21032_/X _26491_/D vssd1 vssd1 vccd1 vccd1 _26491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25442_ _25553_/A vssd1 vssd1 vccd1 vccd1 _25442_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22654_ _22686_/A vssd1 vssd1 vccd1 vccd1 _22654_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21605_ _21599_/X _21600_/X _21601_/X _21602_/X _21603_/X _21604_/X vssd1 vssd1 vccd1
+ vccd1 _21606_/A sky130_fd_sc_hd__mux4_1
XFILLER_159_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22585_ _22577_/X _22578_/X _22579_/X _22580_/X _22581_/X _22582_/X vssd1 vssd1 vccd1
+ vccd1 _22586_/A sky130_fd_sc_hd__mux4_1
X_25373_ _25373_/A vssd1 vssd1 vccd1 vccd1 _27726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27112_ _27112_/CLK _27112_/D vssd1 vssd1 vccd1 vccd1 _27112_/Q sky130_fd_sc_hd__dfxtp_1
X_24324_ _27546_/Q _24328_/B vssd1 vssd1 vccd1 vccd1 _24325_/A sky130_fd_sc_hd__and2_1
X_21536_ _21536_/A vssd1 vssd1 vccd1 vccd1 _21536_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27043_ _22952_/X _27043_/D vssd1 vssd1 vccd1 vccd1 _27043_/Q sky130_fd_sc_hd__dfxtp_1
X_21467_ _21459_/X _21460_/X _21461_/X _21462_/X _21463_/X _21464_/X vssd1 vssd1 vccd1
+ vccd1 _21468_/A sky130_fd_sc_hd__mux4_1
X_24255_ _24255_/A _24256_/B vssd1 vssd1 vccd1 vccd1 _27399_/D sky130_fd_sc_hd__nor2_1
XFILLER_193_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23206_ _23252_/S vssd1 vssd1 vccd1 vccd1 _23215_/S sky130_fd_sc_hd__clkbuf_2
X_20418_ _20408_/X _20409_/X _20410_/X _20411_/X _20412_/X _20413_/X vssd1 vssd1 vccd1
+ vccd1 _20419_/A sky130_fd_sc_hd__mux4_1
X_21398_ _21398_/A vssd1 vssd1 vccd1 vccd1 _21398_/X sky130_fd_sc_hd__clkbuf_1
X_24186_ _24186_/A vssd1 vssd1 vccd1 vccd1 _24195_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_190_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23137_ _27109_/Q _17712_/X _23143_/S vssd1 vssd1 vccd1 vccd1 _23138_/A sky130_fd_sc_hd__mux2_1
X_20349_ _20349_/A vssd1 vssd1 vccd1 vccd1 _20349_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23068_ _27079_/Q _17718_/X _23070_/S vssd1 vssd1 vccd1 vccd1 _23069_/A sky130_fd_sc_hd__mux2_1
X_27945_ _27945_/A _15930_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
XFILLER_49_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22019_ _22019_/A vssd1 vssd1 vccd1 vccd1 _22085_/A sky130_fd_sc_hd__clkbuf_2
X_14910_ _14743_/X _26479_/Q _14918_/S vssd1 vssd1 vccd1 vccd1 _14911_/A sky130_fd_sc_hd__mux2_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _15893_/A vssd1 vssd1 vccd1 vccd1 _15890_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26827_ _22208_/X _26827_/D vssd1 vssd1 vccd1 vccd1 _26827_/Q sky130_fd_sc_hd__dfxtp_1
X_14841_ _14841_/A vssd1 vssd1 vccd1 vccd1 _26510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17560_ _17466_/X _25856_/Q _17562_/S vssd1 vssd1 vccd1 vccd1 _17561_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26758_ _21962_/X _26758_/D vssd1 vssd1 vccd1 vccd1 _26758_/Q sky130_fd_sc_hd__dfxtp_1
X_14772_ _16240_/A vssd1 vssd1 vccd1 vccd1 _14772_/X sky130_fd_sc_hd__buf_2
XFILLER_57_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16511_ _16257_/A _16697_/A _16670_/A _16486_/A vssd1 vssd1 vccd1 vccd1 _16512_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13723_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13778_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_25709_ _25709_/A vssd1 vssd1 vccd1 vccd1 _25709_/X sky130_fd_sc_hd__clkbuf_2
X_17491_ _17491_/A vssd1 vssd1 vccd1 vccd1 _25831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26689_ _21720_/X _26689_/D vssd1 vssd1 vccd1 vccd1 _26689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19230_ _19158_/X _19228_/X _19229_/X vssd1 vssd1 vccd1 vccd1 _19230_/X sky130_fd_sc_hd__o21a_1
X_16442_ _16442_/A _16563_/B vssd1 vssd1 vccd1 vccd1 _16442_/Y sky130_fd_sc_hd__nor2_1
X_13654_ _13923_/A _13661_/B vssd1 vssd1 vccd1 vccd1 _13654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19161_ _26951_/Q _26919_/Q _26887_/Q _26855_/Q _19044_/X _19116_/X vssd1 vssd1 vccd1
+ vccd1 _19161_/X sky130_fd_sc_hd__mux4_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _16851_/A _16851_/B _16703_/A vssd1 vssd1 vccd1 vccd1 _16715_/B sky130_fd_sc_hd__or3b_1
XFILLER_169_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13585_ _14813_/B _13762_/B vssd1 vssd1 vccd1 vccd1 _13602_/A sky130_fd_sc_hd__or2_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112_ _18387_/A vssd1 vssd1 vccd1 vccd1 _18112_/X sky130_fd_sc_hd__clkbuf_2
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15324_ _26302_/Q _13408_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15325_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19092_ _27803_/Q _26564_/Q _26436_/Q _26116_/Q _18974_/X _19019_/X vssd1 vssd1 vccd1
+ vccd1 _19092_/X sky130_fd_sc_hd__mux4_2
XFILLER_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18043_ _18043_/A _17935_/X vssd1 vssd1 vccd1 vccd1 _18043_/X sky130_fd_sc_hd__or2b_1
XFILLER_184_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15255_ _15255_/A vssd1 vssd1 vccd1 vccd1 _26333_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ _26726_/Q _14199_/X _14194_/X _14205_/Y vssd1 vssd1 vccd1 vccd1 _26726_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_193_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15186_ _26363_/Q _13417_/X _15188_/S vssd1 vssd1 vccd1 vccd1 _15187_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ _26751_/Q _14130_/X _14133_/X _14136_/Y vssd1 vssd1 vccd1 vccd1 _26751_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_113_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19994_ _20064_/A vssd1 vssd1 vccd1 vccd1 _19994_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14068_ _14333_/A _14070_/B vssd1 vssd1 vccd1 vccd1 _14068_/Y sky130_fd_sc_hd__nor2_1
X_18945_ _18945_/A vssd1 vssd1 vccd1 vccd1 _19438_/A sky130_fd_sc_hd__buf_2
XFILLER_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _13019_/A vssd1 vssd1 vccd1 vccd1 _13108_/A sky130_fd_sc_hd__clkbuf_4
X_18876_ _26940_/Q _26908_/Q _26876_/Q _26844_/Q _18875_/X _18790_/X vssd1 vssd1 vccd1
+ vccd1 _18876_/X sky130_fd_sc_hd__mux4_2
XFILLER_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17827_ _18379_/A vssd1 vssd1 vccd1 vccd1 _17827_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17758_ _25937_/Q _17756_/X _17770_/S vssd1 vssd1 vccd1 vccd1 _17759_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16709_ _16392_/Y _16399_/Y _16707_/Y _16708_/Y vssd1 vssd1 vccd1 vccd1 _16710_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17689_ _27412_/Q vssd1 vssd1 vccd1 vccd1 _17689_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19428_ _19428_/A vssd1 vssd1 vccd1 vccd1 _19534_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19359_ _19356_/X _19357_/X _19468_/S vssd1 vssd1 vccd1 vccd1 _19359_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22370_ _22435_/A vssd1 vssd1 vccd1 vccd1 _22370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21321_ _21579_/A vssd1 vssd1 vccd1 vccd1 _21389_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24040_ _24038_/X _24039_/X _24047_/S vssd1 vssd1 vccd1 vccd1 _24040_/X sky130_fd_sc_hd__mux2_1
X_21252_ _21252_/A vssd1 vssd1 vccd1 vccd1 _21252_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20203_ _20251_/A vssd1 vssd1 vccd1 vccd1 _20203_/X sky130_fd_sc_hd__clkbuf_1
X_27955__441 vssd1 vssd1 vccd1 vccd1 _27955__441/HI _27955_/A sky130_fd_sc_hd__conb_1
X_21183_ _21199_/A vssd1 vssd1 vccd1 vccd1 _21183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20134_ _20150_/A vssd1 vssd1 vccd1 vccd1 _20134_/X sky130_fd_sc_hd__clkbuf_2
X_25991_ _25991_/CLK _25991_/D vssd1 vssd1 vccd1 vccd1 _25991_/Q sky130_fd_sc_hd__dfxtp_1
X_27730_ _27752_/CLK _27730_/D vssd1 vssd1 vccd1 vccd1 _27730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20065_ _20065_/A vssd1 vssd1 vccd1 vccd1 _20065_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24942_ _25580_/A _24941_/C _24941_/A vssd1 vssd1 vccd1 vccd1 _24943_/B sky130_fd_sc_hd__a21oi_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27661_ _27663_/CLK _27661_/D vssd1 vssd1 vccd1 vccd1 _27661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24873_ _27764_/Q _24873_/B vssd1 vssd1 vccd1 vccd1 _24874_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater260 _27608_/CLK vssd1 vssd1 vccd1 vccd1 _27611_/CLK sky130_fd_sc_hd__clkbuf_1
X_26612_ _21454_/X _26612_/D vssd1 vssd1 vccd1 vccd1 _26612_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater271 _27602_/CLK vssd1 vssd1 vccd1 vccd1 _27488_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater282 _27520_/CLK vssd1 vssd1 vccd1 vccd1 _27523_/CLK sky130_fd_sc_hd__clkbuf_1
X_23824_ _23800_/X _23822_/X _23823_/X _23816_/X vssd1 vssd1 vccd1 vccd1 _27277_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater293 _27262_/CLK vssd1 vssd1 vccd1 vccd1 _27261_/CLK sky130_fd_sc_hd__clkbuf_1
X_27592_ _27592_/CLK _27592_/D vssd1 vssd1 vccd1 vccd1 _27592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_305 _18522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_316 _24400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_327 _24925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 _13204_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26543_ _21208_/X _26543_/D vssd1 vssd1 vccd1 vccd1 _26543_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23755_ _24046_/S vssd1 vssd1 vccd1 vccd1 _23796_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 _16099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20967_ _20953_/X _20954_/X _20955_/X _20956_/X _20958_/X _20960_/X vssd1 vssd1 vccd1
+ vccd1 _20968_/A sky130_fd_sc_hd__mux4_1
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22706_ _22706_/A vssd1 vssd1 vccd1 vccd1 _22706_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26474_ _20970_/X _26474_/D vssd1 vssd1 vccd1 vccd1 _26474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23686_ _24893_/A _27248_/Q _23694_/S vssd1 vssd1 vccd1 vccd1 _23687_/A sky130_fd_sc_hd__mux2_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _20898_/A vssd1 vssd1 vccd1 vccd1 _20898_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25425_ _25425_/A vssd1 vssd1 vccd1 vccd1 _27750_/D sky130_fd_sc_hd__clkbuf_1
X_22637_ _22685_/A vssd1 vssd1 vccd1 vccd1 _22637_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25356_ _25356_/A _25356_/B vssd1 vssd1 vccd1 vccd1 _25356_/Y sky130_fd_sc_hd__nand2_1
X_13370_ _13402_/A vssd1 vssd1 vccd1 vccd1 _13383_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22568_ _22568_/A vssd1 vssd1 vccd1 vccd1 _22568_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24307_ _16131_/X _16133_/Y _16134_/X _24217_/A vssd1 vssd1 vccd1 vccd1 _27436_/D
+ sky130_fd_sc_hd__a31oi_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21519_ _21513_/X _21514_/X _21515_/X _21516_/X _21517_/X _21518_/X vssd1 vssd1 vccd1
+ vccd1 _21520_/A sky130_fd_sc_hd__mux4_1
XFILLER_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25287_ _25287_/A _25287_/B vssd1 vssd1 vccd1 vccd1 _25299_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22499_ _22487_/X _22488_/X _22489_/X _22490_/X _22491_/X _22492_/X vssd1 vssd1 vccd1
+ vccd1 _22500_/A sky130_fd_sc_hd__mux4_1
XFILLER_10_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15040_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27026_ _22900_/X _27026_/D vssd1 vssd1 vccd1 vccd1 _27026_/Q sky130_fd_sc_hd__dfxtp_1
X_24238_ _24238_/A vssd1 vssd1 vccd1 vccd1 _24330_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_170_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24169_ _27461_/Q _24173_/B vssd1 vssd1 vccd1 vccd1 _24170_/A sky130_fd_sc_hd__and2_1
XFILLER_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16991_ input36/X vssd1 vssd1 vccd1 vccd1 _17338_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18730_ _18730_/A vssd1 vssd1 vccd1 vccd1 _26026_/D sky130_fd_sc_hd__clkbuf_1
X_15942_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15942_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_685 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27928_ _27928_/A _15958_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18661_ _25996_/Q _17734_/X _18663_/S vssd1 vssd1 vccd1 vccd1 _18662_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15873_/Y sky130_fd_sc_hd__inv_2
X_27859_ _25810_/X _27859_/D vssd1 vssd1 vccd1 vccd1 _27859_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _26517_/Q _13334_/X _14824_/S vssd1 vssd1 vccd1 vccd1 _14825_/A sky130_fd_sc_hd__mux2_1
X_17612_ _17437_/X _25879_/Q _17612_/S vssd1 vssd1 vccd1 vccd1 _17613_/A sky130_fd_sc_hd__mux2_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18592_ _25572_/A _25582_/A _25583_/A _25584_/A vssd1 vssd1 vccd1 vccd1 _25437_/A
+ sky130_fd_sc_hd__o31ai_2
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17543_ _17440_/X _25848_/Q _17551_/S vssd1 vssd1 vccd1 vccd1 _17544_/A sky130_fd_sc_hd__mux2_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _14755_/A vssd1 vssd1 vccd1 vccd1 _26540_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13706_ _13887_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13706_/Y sky130_fd_sc_hd__nor2_1
X_17474_ _17472_/X _25826_/Q _17486_/S vssd1 vssd1 vccd1 vccd1 _17475_/A sky130_fd_sc_hd__mux2_1
X_14686_ _15758_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_189_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19213_ _26409_/Q _26377_/Q _26345_/Q _26313_/Q _18900_/X _18920_/X vssd1 vssd1 vccd1
+ vccd1 _19213_/X sky130_fd_sc_hd__mux4_1
X_16425_ _16772_/B _16479_/B vssd1 vssd1 vccd1 vccd1 _16890_/B sky130_fd_sc_hd__xnor2_1
X_13637_ _13908_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19144_ _19441_/A vssd1 vssd1 vccd1 vccd1 _19144_/X sky130_fd_sc_hd__buf_2
XFILLER_73_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16356_ _16764_/B vssd1 vssd1 vccd1 vccd1 _16395_/A sky130_fd_sc_hd__clkbuf_1
X_13568_ _14521_/A vssd1 vssd1 vccd1 vccd1 _13934_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_158_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15307_ _15307_/A vssd1 vssd1 vccd1 vccd1 _26310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19075_ _26275_/Q _26243_/Q _26211_/Q _26179_/Q _19028_/X _19074_/X vssd1 vssd1 vccd1
+ vccd1 _19075_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16287_ _16287_/A _16296_/B _26063_/Q vssd1 vssd1 vccd1 vccd1 _16287_/X sky130_fd_sc_hd__or3b_2
X_13499_ _13895_/A _13517_/B vssd1 vssd1 vccd1 vccd1 _13499_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18026_ _18285_/A vssd1 vssd1 vccd1 vccd1 _18026_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15238_ _15238_/A vssd1 vssd1 vccd1 vccd1 _26341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_523 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15169_ _26371_/Q _13392_/X _15173_/S vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_409 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19977_ _19977_/A vssd1 vssd1 vccd1 vccd1 _19977_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18928_ _19555_/A _18928_/B vssd1 vssd1 vccd1 vccd1 _18928_/X sky130_fd_sc_hd__or2_1
XFILLER_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18859_ _19317_/A vssd1 vssd1 vccd1 vccd1 _18859_/X sky130_fd_sc_hd__buf_2
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21870_ _21870_/A vssd1 vssd1 vccd1 vccd1 _21870_/X sky130_fd_sc_hd__clkbuf_1
X_20821_ _20853_/A vssd1 vssd1 vccd1 vccd1 _20821_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23540_ _23543_/A _23540_/B vssd1 vssd1 vccd1 vccd1 _23541_/A sky130_fd_sc_hd__and2_1
X_20752_ _20738_/X _20739_/X _20740_/X _20741_/X _20742_/X _20743_/X vssd1 vssd1 vccd1
+ vccd1 _20753_/A sky130_fd_sc_hd__mux4_1
XFILLER_165_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23471_ input19/X _23469_/X _23470_/X _23461_/X vssd1 vssd1 vccd1 vccd1 _27181_/D
+ sky130_fd_sc_hd__o211a_1
X_20683_ _20683_/A vssd1 vssd1 vccd1 vccd1 _20683_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25210_ _27532_/Q _27500_/Q vssd1 vssd1 vccd1 vccd1 _25211_/B sky130_fd_sc_hd__or2_1
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22422_ _22422_/A vssd1 vssd1 vccd1 vccd1 _22422_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26190_ _19979_/X _26190_/D vssd1 vssd1 vccd1 vccd1 _26190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25141_ _25143_/A vssd1 vssd1 vccd1 vccd1 _25308_/A sky130_fd_sc_hd__clkbuf_2
X_22353_ _22525_/A vssd1 vssd1 vccd1 vccd1 _22422_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21304_ _21304_/A vssd1 vssd1 vccd1 vccd1 _21304_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22284_ _22349_/A vssd1 vssd1 vccd1 vccd1 _22284_/X sky130_fd_sc_hd__clkbuf_1
X_25072_ _25069_/X _25071_/X _25087_/S vssd1 vssd1 vccd1 vccd1 _25072_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24023_ _25940_/Q _26006_/Q _25839_/Q _26038_/Q _23993_/X _23744_/A vssd1 vssd1 vccd1
+ vccd1 _24023_/X sky130_fd_sc_hd__mux4_1
X_21235_ _22543_/A vssd1 vssd1 vccd1 vccd1 _21583_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21166_ _21214_/A vssd1 vssd1 vccd1 vccd1 _21166_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20117_ _20165_/A vssd1 vssd1 vccd1 vccd1 _20117_/X sky130_fd_sc_hd__clkbuf_1
X_25974_ _25974_/CLK _25974_/D vssd1 vssd1 vccd1 vccd1 _25974_/Q sky130_fd_sc_hd__dfxtp_1
X_21097_ _21113_/A vssd1 vssd1 vccd1 vccd1 _21097_/X sky130_fd_sc_hd__clkbuf_2
X_27713_ _27773_/CLK _27713_/D vssd1 vssd1 vccd1 vccd1 _27713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20048_ _20064_/A vssd1 vssd1 vccd1 vccd1 _20048_/X sky130_fd_sc_hd__clkbuf_2
X_24925_ _24925_/A _24925_/B _24925_/C vssd1 vssd1 vccd1 vccd1 _24931_/B sky130_fd_sc_hd__and3_1
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27644_ _27645_/CLK _27644_/D vssd1 vssd1 vccd1 vccd1 _27644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24856_ _27761_/Q _24857_/B vssd1 vssd1 vccd1 vccd1 _24867_/C sky130_fd_sc_hd__and2_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _19345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _22537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23807_ _23803_/X _23805_/X _23844_/S vssd1 vssd1 vccd1 vccd1 _23807_/X sky130_fd_sc_hd__mux2_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _22546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27575_ _27575_/CLK _27575_/D vssd1 vssd1 vccd1 vccd1 _27575_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24787_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24787_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_135 _25810_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21999_ _21999_/A vssd1 vssd1 vccd1 vccd1 _21999_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_146 _13105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _13376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _15701_/A _14542_/B vssd1 vssd1 vccd1 vccd1 _14540_/Y sky130_fd_sc_hd__nor2_1
X_26526_ _21156_/X _26526_/D vssd1 vssd1 vccd1 vccd1 _26526_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _13414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23738_ _27383_/Q _27382_/Q _24061_/A _23035_/C vssd1 vssd1 vccd1 vccd1 _23990_/A
+ sky130_fd_sc_hd__or4b_4
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_179 _16536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14471_ _14471_/A vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__buf_2
X_26457_ _20916_/X _26457_/D vssd1 vssd1 vccd1 vccd1 _26457_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23669_ _23669_/A vssd1 vssd1 vccd1 vccd1 _27240_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16210_ _27382_/Q vssd1 vssd1 vccd1 vccd1 _17420_/B sky130_fd_sc_hd__inv_2
X_25408_ _25408_/A vssd1 vssd1 vccd1 vccd1 _27742_/D sky130_fd_sc_hd__clkbuf_1
X_13422_ _13422_/A vssd1 vssd1 vccd1 vccd1 _26970_/D sky130_fd_sc_hd__clkbuf_1
X_17190_ _17190_/A vssd1 vssd1 vccd1 vccd1 _27930_/A sky130_fd_sc_hd__clkbuf_2
X_26388_ _20665_/X _26388_/D vssd1 vssd1 vccd1 vccd1 _26388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _16151_/A _24306_/A _16845_/A vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__o21ai_1
XFILLER_10_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25339_ _25339_/A _25339_/B vssd1 vssd1 vccd1 vccd1 _25343_/A sky130_fd_sc_hd__nand2_1
X_13353_ _14743_/A vssd1 vssd1 vccd1 vccd1 _13353_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ _16033_/A _16536_/B _16067_/X _16068_/Y _16071_/Y vssd1 vssd1 vccd1 vccd1
+ _16073_/C sky130_fd_sc_hd__o221a_2
XFILLER_6_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13284_ _13284_/A vssd1 vssd1 vccd1 vccd1 _27018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15023_ _15023_/A vssd1 vssd1 vccd1 vccd1 _15034_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19900_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19900_/X sky130_fd_sc_hd__clkbuf_1
X_27009_ _22836_/X _27009_/D vssd1 vssd1 vccd1 vccd1 _27009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19831_ _19898_/A vssd1 vssd1 vccd1 vccd1 _19831_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19762_ _19745_/X _19747_/X _19749_/X _19751_/X _19752_/X _19753_/X vssd1 vssd1 vccd1
+ vccd1 _19763_/A sky130_fd_sc_hd__mux4_1
XFILLER_96_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16974_ _16974_/A vssd1 vssd1 vccd1 vccd1 _16974_/Y sky130_fd_sc_hd__inv_2
X_18713_ _26019_/Q _17705_/X _18713_/S vssd1 vssd1 vccd1 vccd1 _18714_/A sky130_fd_sc_hd__mux2_1
X_15925_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15930_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19693_ _19693_/A vssd1 vssd1 vccd1 vccd1 _19693_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 io_in[9] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18644_ _25988_/Q _17708_/X _18652_/S vssd1 vssd1 vccd1 vccd1 _18645_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15856_ _15980_/A vssd1 vssd1 vccd1 vccd1 _15988_/A sky130_fd_sc_hd__clkbuf_4
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ _14807_/A vssd1 vssd1 vccd1 vccd1 _14807_/X sky130_fd_sc_hd__buf_2
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15787_ _15787_/A vssd1 vssd1 vccd1 vccd1 _26105_/D sky130_fd_sc_hd__clkbuf_1
X_18575_ _18575_/A _18479_/X vssd1 vssd1 vccd1 vccd1 _18575_/X sky130_fd_sc_hd__or2b_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _12999_/A vssd1 vssd1 vccd1 vccd1 _27799_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17526_ _27380_/Q _17674_/C vssd1 vssd1 vccd1 vccd1 _25735_/C sky130_fd_sc_hd__or2_1
X_14738_ _14737_/X _26545_/Q _14741_/S vssd1 vssd1 vccd1 vccd1 _14739_/A sky130_fd_sc_hd__mux2_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17457_ _17524_/S vssd1 vssd1 vccd1 vccd1 _17470_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ _15743_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14669_/Y sky130_fd_sc_hd__nor2_1
X_16408_ _16408_/A vssd1 vssd1 vccd1 vccd1 _16733_/B sky130_fd_sc_hd__clkbuf_2
X_17388_ _17388_/A vssd1 vssd1 vccd1 vccd1 _27947_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19127_ _26533_/Q _26501_/Q _26469_/Q _27045_/Q _19102_/X _19032_/X vssd1 vssd1 vccd1
+ vccd1 _19127_/X sky130_fd_sc_hd__mux4_1
X_16339_ _27376_/Q _16402_/A vssd1 vssd1 vccd1 vccd1 _16339_/X sky130_fd_sc_hd__and2_1
XFILLER_118_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19058_ _19051_/X _19053_/X _19057_/X _19035_/X _18987_/X vssd1 vssd1 vccd1 vccd1
+ _19059_/C sky130_fd_sc_hd__a221o_1
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18009_ _18379_/A vssd1 vssd1 vccd1 vccd1 _18009_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21020_ _21020_/A vssd1 vssd1 vccd1 vccd1 _21020_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22971_ _22955_/X _22956_/X _22957_/X _22958_/X _22960_/X _22962_/X vssd1 vssd1 vccd1
+ vccd1 _22972_/A sky130_fd_sc_hd__mux4_1
XFILLER_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24710_ _24405_/A _24700_/X _24709_/X _24703_/X vssd1 vssd1 vccd1 vccd1 _27601_/D
+ sky130_fd_sc_hd__o211a_1
X_21922_ _21922_/A vssd1 vssd1 vccd1 vccd1 _21922_/X sky130_fd_sc_hd__clkbuf_1
X_25690_ _25722_/A vssd1 vssd1 vccd1 vccd1 _25690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24641_ _24748_/A vssd1 vssd1 vccd1 vccd1 _24841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21853_ _21844_/X _21846_/X _21848_/X _21850_/X _21851_/X _21852_/X vssd1 vssd1 vccd1
+ vccd1 _21854_/A sky130_fd_sc_hd__mux4_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20804_ _20852_/A vssd1 vssd1 vccd1 vccd1 _20804_/X sky130_fd_sc_hd__clkbuf_2
X_27360_ _27478_/CLK _27360_/D vssd1 vssd1 vccd1 vccd1 _27360_/Q sky130_fd_sc_hd__dfxtp_1
X_24572_ _27647_/Q _24576_/B vssd1 vssd1 vccd1 vccd1 _24573_/A sky130_fd_sc_hd__and2_1
X_21784_ _21784_/A vssd1 vssd1 vccd1 vccd1 _21784_/X sky130_fd_sc_hd__clkbuf_1
X_26311_ _20401_/X _26311_/D vssd1 vssd1 vccd1 vccd1 _26311_/Q sky130_fd_sc_hd__dfxtp_1
X_23523_ _23523_/A vssd1 vssd1 vccd1 vccd1 _27198_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27291_ _27299_/CLK _27291_/D vssd1 vssd1 vccd1 vccd1 _27291_/Q sky130_fd_sc_hd__dfxtp_1
X_20735_ _20735_/A vssd1 vssd1 vccd1 vccd1 _20735_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26242_ _20157_/X _26242_/D vssd1 vssd1 vccd1 vccd1 _26242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23454_ input13/X _23442_/X _23453_/X _23447_/X vssd1 vssd1 vccd1 vccd1 _27175_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20666_ _20652_/X _20653_/X _20654_/X _20655_/X _20656_/X _20657_/X vssd1 vssd1 vccd1
+ vccd1 _20667_/A sky130_fd_sc_hd__mux4_1
XFILLER_177_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22405_ _22421_/A vssd1 vssd1 vccd1 vccd1 _22405_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26173_ _19913_/X _26173_/D vssd1 vssd1 vccd1 vccd1 _26173_/Q sky130_fd_sc_hd__dfxtp_1
X_23385_ _24767_/A _27246_/Q _27235_/Q _24733_/A vssd1 vssd1 vccd1 vccd1 _23385_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_20597_ _20597_/A vssd1 vssd1 vccd1 vccd1 _20597_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25124_ _27691_/Q _25112_/X _25123_/Y _23498_/X vssd1 vssd1 vccd1 vccd1 _27691_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_192_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22336_ _22336_/A vssd1 vssd1 vccd1 vccd1 _22336_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25055_ _25051_/X _25053_/X _25087_/S vssd1 vssd1 vccd1 vccd1 _25055_/X sky130_fd_sc_hd__mux2_1
X_22267_ _22525_/A vssd1 vssd1 vccd1 vccd1 _22336_/A sky130_fd_sc_hd__clkbuf_2
X_24006_ _23990_/X _24000_/X _24004_/X _24005_/X vssd1 vssd1 vccd1 vccd1 _27296_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21218_ _21290_/A vssd1 vssd1 vccd1 vccd1 _21218_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22198_ _22263_/A vssd1 vssd1 vccd1 vccd1 _22198_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21149_ _21149_/A vssd1 vssd1 vccd1 vccd1 _21214_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _14348_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _13971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25957_ _27325_/CLK _25957_/D vssd1 vssd1 vccd1 vccd1 _25957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15710_ _15710_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15710_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12922_ input41/X input52/X input63/X input66/X vssd1 vssd1 vccd1 vccd1 _23325_/A
+ sky130_fd_sc_hd__or4_1
X_24908_ _27658_/Q _24885_/X _24907_/Y _24890_/X vssd1 vssd1 vccd1 vccd1 _27658_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16690_ _16779_/A _16688_/Y _16689_/X vssd1 vssd1 vccd1 vccd1 _16690_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25888_ _25925_/CLK _25888_/D vssd1 vssd1 vccd1 vccd1 _25888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15641_ _13099_/X _26162_/Q _15645_/S vssd1 vssd1 vccd1 vccd1 _15642_/A sky130_fd_sc_hd__mux2_1
X_27627_ _27627_/CLK _27627_/D vssd1 vssd1 vccd1 vccd1 _27627_/Q sky130_fd_sc_hd__dfxtp_1
X_24839_ _24914_/A vssd1 vssd1 vccd1 vccd1 _24839_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18360_/A vssd1 vssd1 vccd1 vccd1 _18360_/X sky130_fd_sc_hd__buf_2
XFILLER_15_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27558_ _27558_/CLK _27558_/D vssd1 vssd1 vccd1 vccd1 _27558_/Q sky130_fd_sc_hd__dfxtp_1
X_15572_ _15572_/A vssd1 vssd1 vccd1 vccd1 _26193_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17311_ _27219_/Q _17310_/X _17311_/S vssd1 vssd1 vccd1 vccd1 _17312_/A sky130_fd_sc_hd__mux2_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _26621_/Q _14514_/X _14510_/X _14522_/Y vssd1 vssd1 vccd1 vccd1 _26621_/D
+ sky130_fd_sc_hd__a31o_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26509_ _21092_/X _26509_/D vssd1 vssd1 vccd1 vccd1 _26509_/Q sky130_fd_sc_hd__dfxtp_1
X_18291_ _18289_/X _18290_/X _18514_/S vssd1 vssd1 vccd1 vccd1 _18291_/X sky130_fd_sc_hd__mux2_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27489_ _27534_/CLK _27489_/D vssd1 vssd1 vccd1 vccd1 _27489_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17303_/A vssd1 vssd1 vccd1 vccd1 _17242_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14454_ _26640_/Q _14441_/X _14437_/X _14453_/Y vssd1 vssd1 vccd1 vccd1 _26640_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13405_ _16224_/A vssd1 vssd1 vccd1 vccd1 _13405_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_179_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17173_ _27079_/Q _27111_/Q _17173_/S vssd1 vssd1 vccd1 vccd1 _17173_/X sky130_fd_sc_hd__mux2_1
X_14385_ _14398_/A vssd1 vssd1 vccd1 vccd1 _14385_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16124_ _16151_/A _24309_/A vssd1 vssd1 vccd1 vccd1 _16125_/B sky130_fd_sc_hd__or2_1
XFILLER_116_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_592 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13336_ _13336_/A vssd1 vssd1 vccd1 vccd1 _26997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16055_ _16047_/Y _13672_/A _16054_/X vssd1 vssd1 vccd1 vccd1 _16313_/B sky130_fd_sc_hd__o21ba_1
X_13267_ _27025_/Q _13105_/X _13269_/S vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15006_ _15743_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _16206_/A vssd1 vssd1 vccd1 vccd1 _13198_/X sky130_fd_sc_hd__buf_2
XFILLER_155_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19814_ _19814_/A vssd1 vssd1 vccd1 vccd1 _19814_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19745_ _19812_/A vssd1 vssd1 vccd1 vccd1 _19745_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16957_ _24635_/A _24488_/B vssd1 vssd1 vccd1 vccd1 _24522_/A sky130_fd_sc_hd__and2_1
XFILLER_38_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15908_ _15912_/A vssd1 vssd1 vccd1 vccd1 _15908_/Y sky130_fd_sc_hd__inv_2
X_19676_ _19659_/X _19661_/X _19663_/X _19665_/X _19666_/X _19667_/X vssd1 vssd1 vccd1
+ vccd1 _19677_/A sky130_fd_sc_hd__mux4_1
X_16888_ _16888_/A _16888_/B vssd1 vssd1 vccd1 vccd1 _16888_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18627_ _18627_/A vssd1 vssd1 vccd1 vccd1 _25980_/D sky130_fd_sc_hd__clkbuf_1
X_15839_ _15839_/A vssd1 vssd1 vccd1 vccd1 _26081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18558_ _26296_/Q _26264_/Q _26232_/Q _26200_/Q _18458_/X _18481_/X vssd1 vssd1 vccd1
+ vccd1 _18558_/X sky130_fd_sc_hd__mux4_1
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17509_ _17508_/X _25837_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17510_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18489_ _18489_/A vssd1 vssd1 vccd1 vccd1 _18489_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_13 _25925_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20520_ _20512_/X _20513_/X _20514_/X _20515_/X _20517_/X _20519_/X vssd1 vssd1 vccd1
+ vccd1 _20521_/A sky130_fd_sc_hd__mux4_1
XANTENNA_24 _27141_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_35 _18458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 _17952_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_57 _18224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20451_ _20515_/A vssd1 vssd1 vccd1 vccd1 _20451_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_68 _18340_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_79 _18782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23170_ _27124_/Q _17760_/X _23176_/S vssd1 vssd1 vccd1 vccd1 _23171_/A sky130_fd_sc_hd__mux2_1
X_20382_ _20376_/X _20377_/X _20378_/X _20379_/X _20380_/X _20381_/X vssd1 vssd1 vccd1
+ vccd1 _20383_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22121_ _22103_/X _22106_/X _22109_/X _22112_/X _22113_/X _22114_/X vssd1 vssd1 vccd1
+ vccd1 _22122_/A sky130_fd_sc_hd__mux4_1
XFILLER_161_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22052_ _22084_/A vssd1 vssd1 vccd1 vccd1 _22052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21003_ _20991_/X _20992_/X _20993_/X _20994_/X _20995_/X _20996_/X vssd1 vssd1 vccd1
+ vccd1 _21004_/A sky130_fd_sc_hd__mux4_1
XFILLER_88_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26860_ _22322_/X _26860_/D vssd1 vssd1 vccd1 vccd1 _26860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25811_ _27129_/CLK _25811_/D vssd1 vssd1 vccd1 vccd1 _25811_/Q sky130_fd_sc_hd__dfxtp_1
X_26791_ _22076_/X _26791_/D vssd1 vssd1 vccd1 vccd1 _26791_/Q sky130_fd_sc_hd__dfxtp_1
X_25742_ _17431_/X _27828_/Q _25746_/S vssd1 vssd1 vccd1 vccd1 _25743_/A sky130_fd_sc_hd__mux2_1
X_22954_ _22954_/A vssd1 vssd1 vccd1 vccd1 _22954_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21905_ _21895_/X _21896_/X _21897_/X _21898_/X _21899_/X _21900_/X vssd1 vssd1 vccd1
+ vccd1 _21906_/A sky130_fd_sc_hd__mux4_1
X_25673_ _25721_/A vssd1 vssd1 vccd1 vccd1 _25673_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22885_ _22869_/X _22870_/X _22871_/X _22872_/X _22874_/X _22876_/X vssd1 vssd1 vccd1
+ vccd1 _22886_/A sky130_fd_sc_hd__mux4_1
XFILLER_83_584 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27412_ _27412_/CLK _27412_/D vssd1 vssd1 vccd1 vccd1 _27412_/Q sky130_fd_sc_hd__dfxtp_1
X_24624_ _27671_/Q _24624_/B vssd1 vssd1 vccd1 vccd1 _24625_/A sky130_fd_sc_hd__and2_1
X_21836_ _21836_/A vssd1 vssd1 vccd1 vccd1 _21836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27343_ _27447_/CLK _27343_/D vssd1 vssd1 vccd1 vccd1 _27343_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24555_ _24555_/A vssd1 vssd1 vccd1 vccd1 _27539_/D sky130_fd_sc_hd__clkbuf_1
X_21767_ _21758_/X _21760_/X _21762_/X _21764_/X _21765_/X _21766_/X vssd1 vssd1 vccd1
+ vccd1 _21768_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23506_ _23562_/A vssd1 vssd1 vccd1 vccd1 _23526_/A sky130_fd_sc_hd__clkbuf_1
X_20718_ _20703_/X _20705_/X _20707_/X _20709_/X _20710_/X _20711_/X vssd1 vssd1 vccd1
+ vccd1 _20719_/A sky130_fd_sc_hd__mux4_1
X_27274_ _27278_/CLK _27274_/D vssd1 vssd1 vccd1 vccd1 _27274_/Q sky130_fd_sc_hd__dfxtp_1
X_24486_ _24486_/A vssd1 vssd1 vccd1 vccd1 _27518_/D sky130_fd_sc_hd__clkbuf_1
X_21698_ _21698_/A vssd1 vssd1 vccd1 vccd1 _21698_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26225_ _20105_/X _26225_/D vssd1 vssd1 vccd1 vccd1 _26225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23437_ _16985_/X _23429_/X _23436_/X _23434_/X vssd1 vssd1 vccd1 vccd1 _27168_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_184_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20649_ _20649_/A vssd1 vssd1 vccd1 vccd1 _20649_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14170_ _14348_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26156_ _19859_/X _26156_/D vssd1 vssd1 vccd1 vccd1 _26156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23368_ _24906_/A _23365_/Y _27260_/Q _24806_/A _23367_/X vssd1 vssd1 vccd1 vccd1
+ _23368_/X sky130_fd_sc_hd__a221o_1
XFILLER_192_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25107_ _25107_/A vssd1 vssd1 vccd1 vccd1 _27753_/D sky130_fd_sc_hd__clkbuf_1
X_13121_ _27355_/Q _13090_/X _13091_/X _27323_/Q _13120_/X vssd1 vssd1 vccd1 vccd1
+ _14747_/A sky130_fd_sc_hd__a221o_4
X_22319_ _22335_/A vssd1 vssd1 vccd1 vccd1 _22319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26087_ _19616_/X _26087_/D vssd1 vssd1 vccd1 vccd1 _26087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23299_ _27736_/Q _23295_/Y _23291_/Y input49/X vssd1 vssd1 vccd1 vccd1 _23299_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13052_ _27065_/Q _13038_/X _13079_/S vssd1 vssd1 vccd1 vccd1 _13053_/A sky130_fd_sc_hd__mux2_1
X_25038_ _25036_/X _25037_/X _25046_/S vssd1 vssd1 vccd1 vccd1 _25038_/X sky130_fd_sc_hd__mux2_1
X_17860_ _27794_/Q _26555_/Q _26427_/Q _26107_/Q _17782_/X _17785_/X vssd1 vssd1 vccd1
+ vccd1 _17860_/X sky130_fd_sc_hd__mux4_2
XFILLER_120_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16811_ _16806_/X _16807_/Y _16811_/C _16811_/D vssd1 vssd1 vccd1 vccd1 _16812_/B
+ sky130_fd_sc_hd__and4bb_1
X_17791_ _18425_/A vssd1 vssd1 vccd1 vccd1 _17791_/X sky130_fd_sc_hd__buf_2
X_26989_ _22766_/X _26989_/D vssd1 vssd1 vccd1 vccd1 _26989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19530_ _19524_/X _19526_/X _19529_/X _19448_/X _19469_/X vssd1 vssd1 vccd1 vccd1
+ _19531_/C sky130_fd_sc_hd__a221o_1
X_13954_ _14335_/A _13954_/B vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16742_ _16742_/A vssd1 vssd1 vccd1 vccd1 _16743_/B sky130_fd_sc_hd__inv_2
XFILLER_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16673_ _16669_/Y _16670_/Y _16672_/Y _16619_/X vssd1 vssd1 vccd1 vccd1 _24243_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_19461_ _26164_/Q _26100_/Q _27028_/Q _26996_/Q _19460_/X _19348_/X vssd1 vssd1 vccd1
+ vccd1 _19462_/B sky130_fd_sc_hd__mux4_1
X_13885_ _26832_/Q _13880_/X _13873_/X _13884_/Y vssd1 vssd1 vccd1 vccd1 _26832_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18412_ _18412_/A vssd1 vssd1 vccd1 vccd1 _18412_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _15680_/A vssd1 vssd1 vccd1 vccd1 _15693_/S sky130_fd_sc_hd__clkbuf_2
X_19392_ _19389_/X _19390_/X _19480_/S vssd1 vssd1 vccd1 vccd1 _19392_/X sky130_fd_sc_hd__mux2_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _26158_/Q _26094_/Q _27022_/Q _26990_/Q _18000_/A _17959_/A vssd1 vssd1 vccd1
+ vccd1 _18344_/A sky130_fd_sc_hd__mux4_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15555_/A vssd1 vssd1 vccd1 vccd1 _26201_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _26626_/Q _14496_/X _14492_/X _14505_/Y vssd1 vssd1 vccd1 vccd1 _26626_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18274_ _18274_/A _18156_/X vssd1 vssd1 vccd1 vccd1 _18274_/X sky130_fd_sc_hd__or2b_1
XFILLER_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15486_ _13067_/X _26231_/Q _15490_/S vssd1 vssd1 vccd1 vccd1 _15487_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14437_ _14510_/A vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17225_ _27212_/Q _17224_/X _17250_/S vssd1 vssd1 vccd1 vccd1 _17226_/A sky130_fd_sc_hd__mux2_1
Xinput11 la1_data_in[11] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput22 la1_data_in[21] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_4
Xinput33 la1_data_in[31] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
X_17156_ _25924_/Q _25990_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17157_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput44 la1_oenb[12] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_8
Xinput55 la1_oenb[22] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_4
X_14368_ _26668_/Q _14365_/X _14358_/X _14367_/Y vssd1 vssd1 vccd1 vccd1 _26668_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 la1_oenb[3] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
X_16107_ _16623_/A vssd1 vssd1 vccd1 vccd1 _16845_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13319_ _14709_/A vssd1 vssd1 vccd1 vccd1 _13319_/X sky130_fd_sc_hd__buf_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17087_ _17057_/X _17086_/X _17033_/X vssd1 vssd1 vccd1 vccd1 _17087_/X sky130_fd_sc_hd__a21bo_1
X_14299_ _26693_/Q _14296_/X _14297_/X _14298_/Y vssd1 vssd1 vccd1 vccd1 _26693_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_196_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16038_ _27478_/Q _27477_/Q vssd1 vssd1 vccd1 vccd1 _16062_/A sky130_fd_sc_hd__or2_1
XFILLER_170_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17989_ _17987_/X _17988_/X _18075_/S vssd1 vssd1 vccd1 vccd1 _17989_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19728_ _19728_/A vssd1 vssd1 vccd1 vccd1 _19728_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19659_ _19726_/A vssd1 vssd1 vccd1 vccd1 _19659_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22670_ _22686_/A vssd1 vssd1 vccd1 vccd1 _22670_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21621_ _21615_/X _21616_/X _21617_/X _21618_/X _21619_/X _21620_/X vssd1 vssd1 vccd1
+ vccd1 _21622_/A sky130_fd_sc_hd__mux4_1
XFILLER_179_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24340_ _24340_/A vssd1 vssd1 vccd1 vccd1 _27453_/D sky130_fd_sc_hd__clkbuf_1
X_21552_ _21552_/A vssd1 vssd1 vccd1 vccd1 _21552_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20503_ _20503_/A vssd1 vssd1 vccd1 vccd1 _20503_/X sky130_fd_sc_hd__clkbuf_1
X_24271_ _16173_/X _16176_/Y _16177_/X _24269_/X vssd1 vssd1 vccd1 vccd1 _27409_/D
+ sky130_fd_sc_hd__o31a_1
X_21483_ _21475_/X _21476_/X _21477_/X _21478_/X _21480_/X _21482_/X vssd1 vssd1 vccd1
+ vccd1 _21484_/A sky130_fd_sc_hd__mux4_1
XFILLER_21_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26010_ _27129_/CLK _26010_/D vssd1 vssd1 vccd1 vccd1 _26010_/Q sky130_fd_sc_hd__dfxtp_1
X_23222_ _17479_/X _27147_/Q _23226_/S vssd1 vssd1 vccd1 vccd1 _23223_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20434_ _20424_/X _20425_/X _20426_/X _20427_/X _20430_/X _20433_/X vssd1 vssd1 vccd1
+ vccd1 _20435_/A sky130_fd_sc_hd__mux4_1
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23153_ _23153_/A vssd1 vssd1 vccd1 vccd1 _27116_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20365_ _20413_/A vssd1 vssd1 vccd1 vccd1 _20365_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22104_ _22540_/A vssd1 vssd1 vccd1 vccd1 _22453_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23084_ _27086_/Q _17740_/X _23092_/S vssd1 vssd1 vccd1 vccd1 _23085_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27961_ _27961_/A _15872_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
X_20296_ _20286_/X _20287_/X _20288_/X _20289_/X _20290_/X _20291_/X vssd1 vssd1 vccd1
+ vccd1 _20297_/A sky130_fd_sc_hd__mux4_1
XFILLER_103_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22035_ _22083_/A vssd1 vssd1 vccd1 vccd1 _22035_/X sky130_fd_sc_hd__clkbuf_1
X_26912_ _22498_/X _26912_/D vssd1 vssd1 vccd1 vccd1 _26912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26843_ _22258_/X _26843_/D vssd1 vssd1 vccd1 vccd1 _26843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26774_ _22014_/X _26774_/D vssd1 vssd1 vccd1 vccd1 _26774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23986_ _27090_/Q _27122_/Q _23986_/S vssd1 vssd1 vccd1 vccd1 _23986_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25725_ _25725_/A vssd1 vssd1 vccd1 vccd1 _25725_/X sky130_fd_sc_hd__clkbuf_2
X_22937_ _22923_/X _22924_/X _22925_/X _22926_/X _22927_/X _22928_/X vssd1 vssd1 vccd1
+ vccd1 _22938_/A sky130_fd_sc_hd__mux4_1
XFILLER_29_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _13940_/A _13670_/B vssd1 vssd1 vccd1 vccd1 _13670_/Y sky130_fd_sc_hd__nor2_1
X_25656_ _25722_/A vssd1 vssd1 vccd1 vccd1 _25656_/X sky130_fd_sc_hd__clkbuf_1
X_22868_ _22868_/A vssd1 vssd1 vccd1 vccd1 _22868_/X sky130_fd_sc_hd__clkbuf_1
X_24607_ _27663_/Q _24609_/B vssd1 vssd1 vccd1 vccd1 _24608_/A sky130_fd_sc_hd__and2_1
X_21819_ _21809_/X _21810_/X _21811_/X _21812_/X _21813_/X _21814_/X vssd1 vssd1 vccd1
+ vccd1 _21820_/A sky130_fd_sc_hd__mux4_1
X_25587_ _27714_/Q _25568_/X _25569_/X vssd1 vssd1 vccd1 vccd1 _25587_/Y sky130_fd_sc_hd__a21oi_1
X_22799_ _22783_/X _22784_/X _22785_/X _22786_/X _22788_/X _22790_/X vssd1 vssd1 vccd1
+ vccd1 _22800_/A sky130_fd_sc_hd__mux4_1
XFILLER_189_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27326_ _27326_/CLK _27326_/D vssd1 vssd1 vccd1 vccd1 _27326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15340_ _14715_/X _26296_/Q _15346_/S vssd1 vssd1 vccd1 vccd1 _15341_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24538_ _24538_/A vssd1 vssd1 vccd1 vccd1 _24552_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27257_ _27783_/CLK _27257_/D vssd1 vssd1 vccd1 vccd1 _27257_/Q sky130_fd_sc_hd__dfxtp_1
X_15271_ _26326_/Q _13331_/X _15273_/S vssd1 vssd1 vccd1 vccd1 _15272_/A sky130_fd_sc_hd__mux2_1
X_24469_ _24480_/A vssd1 vssd1 vccd1 vccd1 _24478_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17010_ _25358_/B vssd1 vssd1 vccd1 vccd1 _17387_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_184_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14222_ _26720_/Q _14212_/X _14220_/X _14221_/Y vssd1 vssd1 vccd1 vccd1 _26720_/D
+ sky130_fd_sc_hd__a31o_1
X_26208_ _20041_/X _26208_/D vssd1 vssd1 vccd1 vccd1 _26208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27188_ _27190_/CLK _27188_/D vssd1 vssd1 vccd1 vccd1 _27188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14153_ _14331_/A _14158_/B vssd1 vssd1 vccd1 vccd1 _14153_/Y sky130_fd_sc_hd__nor2_1
X_26139_ _19795_/X _26139_/D vssd1 vssd1 vccd1 vccd1 _26139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13104_ _27358_/Q _13021_/A _13102_/X _27326_/Q _13103_/X vssd1 vssd1 vccd1 vccd1
+ _14737_/A sky130_fd_sc_hd__a221o_4
X_14084_ _26771_/Q _14076_/X _14080_/X _14083_/Y vssd1 vssd1 vccd1 vccd1 _26771_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18961_ _26526_/Q _26494_/Q _26462_/Q _27038_/Q _18829_/X _18863_/X vssd1 vssd1 vccd1
+ vccd1 _18961_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13169_/B vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__clkbuf_1
X_17912_ _18479_/A vssd1 vssd1 vccd1 vccd1 _17912_/X sky130_fd_sc_hd__clkbuf_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18892_ _18989_/A _18892_/B _18892_/C vssd1 vssd1 vccd1 vccd1 _18893_/A sky130_fd_sc_hd__and3_1
X_17843_ _18141_/A vssd1 vssd1 vccd1 vccd1 _17843_/X sky130_fd_sc_hd__buf_4
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _17774_/A vssd1 vssd1 vccd1 vccd1 _25942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14986_ _15725_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14986_/Y sky130_fd_sc_hd__nor2_1
X_19513_ _19567_/A _19513_/B _19513_/C vssd1 vssd1 vccd1 vccd1 _19514_/A sky130_fd_sc_hd__and3_1
XFILLER_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _24230_/A _24231_/A vssd1 vssd1 vccd1 vccd1 _16874_/C sky130_fd_sc_hd__and2_1
X_13937_ _26812_/Q _13933_/X _13925_/X _13936_/Y vssd1 vssd1 vccd1 vccd1 _26812_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19444_ _26419_/Q _26387_/Q _26355_/Q _26323_/Q _19331_/X _19399_/X vssd1 vssd1 vccd1
+ vccd1 _19444_/X sky130_fd_sc_hd__mux4_1
X_13868_ _13868_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13868_/Y sky130_fd_sc_hd__nor2_1
X_16656_ _24250_/A _24247_/A _24259_/A _24258_/A vssd1 vssd1 vccd1 vccd1 _16896_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_16_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15607_ _15607_/A vssd1 vssd1 vccd1 vccd1 _26177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19375_ _19373_/X _19374_/X _19553_/S vssd1 vssd1 vccd1 vccd1 _19375_/X sky130_fd_sc_hd__mux2_2
X_13799_ _13891_/A _13799_/B vssd1 vssd1 vccd1 vccd1 _13799_/Y sky130_fd_sc_hd__nor2_1
X_16587_ _16888_/A _16571_/X _16573_/X _16586_/X vssd1 vssd1 vccd1 vccd1 _16879_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18326_ _18483_/A vssd1 vssd1 vccd1 vccd1 _18326_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15538_/A vssd1 vssd1 vccd1 vccd1 _26208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18257_ _26282_/Q _26250_/Q _26218_/Q _26186_/Q _18185_/X _18209_/X vssd1 vssd1 vccd1
+ vccd1 _18257_/X sky130_fd_sc_hd__mux4_1
X_15469_ _26238_/Q _13408_/X _15473_/S vssd1 vssd1 vccd1 vccd1 _15470_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17208_ _25827_/Q _26026_/Q _17219_/S vssd1 vssd1 vccd1 vccd1 _17208_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18188_ _26535_/Q _26503_/Q _26471_/Q _27047_/Q _18117_/X _18141_/X vssd1 vssd1 vccd1
+ vccd1 _18188_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17139_ _17387_/S vssd1 vssd1 vccd1 vccd1 _17189_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20150_ _20150_/A vssd1 vssd1 vccd1 vccd1 _20150_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_537 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20081_ _20150_/A vssd1 vssd1 vccd1 vccd1 _20081_/X sky130_fd_sc_hd__clkbuf_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater420 _27331_/CLK vssd1 vssd1 vccd1 vccd1 _27392_/CLK sky130_fd_sc_hd__clkbuf_2
Xrepeater431 _25963_/CLK vssd1 vssd1 vccd1 vccd1 _25969_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23840_ _27074_/Q _23812_/X _23813_/X _27106_/Q _23814_/X vssd1 vssd1 vccd1 vccd1
+ _23840_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27988__454 vssd1 vssd1 vccd1 vccd1 _27988__454/HI _27988_/A sky130_fd_sc_hd__conb_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23771_ _25913_/Q _25979_/Q _25812_/Q _26011_/Q _23747_/X _23749_/X vssd1 vssd1 vccd1
+ vccd1 _23771_/X sky130_fd_sc_hd__mux4_1
X_20983_ _20972_/X _20974_/X _20976_/X _20978_/X _20979_/X _20980_/X vssd1 vssd1 vccd1
+ vccd1 _20984_/A sky130_fd_sc_hd__mux4_1
XFILLER_129_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25510_ _25569_/A vssd1 vssd1 vccd1 vccd1 _25510_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22722_ _22786_/A vssd1 vssd1 vccd1 vccd1 _22722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26490_ _21030_/X _26490_/D vssd1 vssd1 vccd1 vccd1 _26490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25441_ _25583_/A vssd1 vssd1 vccd1 vccd1 _25553_/A sky130_fd_sc_hd__clkbuf_1
X_22653_ _22685_/A vssd1 vssd1 vccd1 vccd1 _22653_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21604_ _21636_/A vssd1 vssd1 vccd1 vccd1 _21604_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25372_ _27726_/Q input68/X _25380_/S vssd1 vssd1 vccd1 vccd1 _25373_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22584_ _22584_/A vssd1 vssd1 vccd1 vccd1 _22584_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27111_ _27111_/CLK _27111_/D vssd1 vssd1 vccd1 vccd1 _27111_/Q sky130_fd_sc_hd__dfxtp_1
X_24323_ _24323_/A vssd1 vssd1 vccd1 vccd1 _27445_/D sky130_fd_sc_hd__clkbuf_1
X_21535_ _21529_/X _21530_/X _21531_/X _21532_/X _21533_/X _21534_/X vssd1 vssd1 vccd1
+ vccd1 _21536_/A sky130_fd_sc_hd__mux4_1
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27042_ _22950_/X _27042_/D vssd1 vssd1 vccd1 vccd1 _27042_/Q sky130_fd_sc_hd__dfxtp_1
X_24254_ _24254_/A vssd1 vssd1 vccd1 vccd1 _27398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21466_ _21466_/A vssd1 vssd1 vccd1 vccd1 _21466_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23205_ _23205_/A vssd1 vssd1 vccd1 vccd1 _27139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20417_ _20417_/A vssd1 vssd1 vccd1 vccd1 _20417_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24185_ _24185_/A vssd1 vssd1 vccd1 vccd1 _27363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21397_ _21389_/X _21390_/X _21391_/X _21392_/X _21394_/X _21396_/X vssd1 vssd1 vccd1
+ vccd1 _21398_/A sky130_fd_sc_hd__mux4_1
XFILLER_190_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23136_ _23136_/A vssd1 vssd1 vccd1 vccd1 _27108_/D sky130_fd_sc_hd__clkbuf_1
X_20348_ _20334_/X _20335_/X _20336_/X _20337_/X _20339_/X _20341_/X vssd1 vssd1 vccd1
+ vccd1 _20349_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_812 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23067_ _23067_/A vssd1 vssd1 vccd1 vccd1 _27078_/D sky130_fd_sc_hd__clkbuf_1
X_27944_ _27944_/A _15933_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
X_20279_ _20279_/A vssd1 vssd1 vccd1 vccd1 _20279_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22018_ _22084_/A vssd1 vssd1 vccd1 vccd1 _22018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26826_ _22206_/X _26826_/D vssd1 vssd1 vccd1 vccd1 _26826_/Q sky130_fd_sc_hd__dfxtp_1
X_14840_ _26510_/Q _13357_/X _14846_/S vssd1 vssd1 vccd1 vccd1 _14841_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14771_ _14771_/A vssd1 vssd1 vccd1 vccd1 _26535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26757_ _21960_/X _26757_/D vssd1 vssd1 vccd1 vccd1 _26757_/Q sky130_fd_sc_hd__dfxtp_1
X_23969_ _25934_/Q _26000_/Q _25833_/Q _26032_/Q _23946_/X _23929_/X vssd1 vssd1 vccd1
+ vccd1 _23969_/X sky130_fd_sc_hd__mux4_1
X_13722_ _26889_/Q _13710_/X _13718_/X _13721_/Y vssd1 vssd1 vccd1 vccd1 _26889_/D
+ sky130_fd_sc_hd__a31o_1
X_16510_ _16666_/B vssd1 vssd1 vccd1 vccd1 _16816_/B sky130_fd_sc_hd__inv_2
XFILLER_72_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25708_ _25724_/A vssd1 vssd1 vccd1 vccd1 _25708_/X sky130_fd_sc_hd__clkbuf_1
X_17490_ _17488_/X _25831_/Q _17502_/S vssd1 vssd1 vccd1 vccd1 _17491_/A sky130_fd_sc_hd__mux2_1
X_26688_ _21718_/X _26688_/D vssd1 vssd1 vccd1 vccd1 _26688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13653_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13653_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16441_ _16779_/B _16441_/B vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__xnor2_1
X_25639_ _25639_/A vssd1 vssd1 vccd1 vccd1 _25709_/A sky130_fd_sc_hd__clkbuf_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19160_ _19158_/X _19159_/X _19089_/X vssd1 vssd1 vccd1 vccd1 _19160_/X sky130_fd_sc_hd__o21a_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16372_/A _16396_/B vssd1 vssd1 vccd1 vccd1 _16703_/A sky130_fd_sc_hd__xnor2_1
X_13584_ _26938_/Q _13580_/X _13442_/B _13583_/Y vssd1 vssd1 vccd1 vccd1 _26938_/D
+ sky130_fd_sc_hd__a31o_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _17972_/X _18104_/X _18109_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _18124_/B
+ sky130_fd_sc_hd__a211o_1
X_15323_ _15323_/A vssd1 vssd1 vccd1 vccd1 _26303_/D sky130_fd_sc_hd__clkbuf_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27309_ _27311_/CLK _27309_/D vssd1 vssd1 vccd1 vccd1 _27309_/Q sky130_fd_sc_hd__dfxtp_1
X_19091_ _26948_/Q _26916_/Q _26884_/Q _26852_/Q _19044_/X _18972_/X vssd1 vssd1 vccd1
+ vccd1 _19091_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15254_ _14801_/X _26333_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15255_/A sky130_fd_sc_hd__mux2_1
X_18042_ _26145_/Q _26081_/Q _27009_/Q _26977_/Q _18041_/X _17959_/X vssd1 vssd1 vccd1
+ vccd1 _18043_/A sky130_fd_sc_hd__mux4_1
XFILLER_200_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14205_ _14383_/A _14213_/B vssd1 vssd1 vccd1 vccd1 _14205_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15185_ _15185_/A vssd1 vssd1 vccd1 vccd1 _26364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _14401_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19993_ _20338_/A vssd1 vssd1 vccd1 vccd1 _20064_/A sky130_fd_sc_hd__buf_2
XFILLER_67_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _26777_/Q _14058_/X _14064_/X _14066_/Y vssd1 vssd1 vccd1 vccd1 _26777_/D
+ sky130_fd_sc_hd__a31o_1
X_18944_ _27797_/Q _26558_/Q _26430_/Q _26110_/Q _18793_/X _18851_/X vssd1 vssd1 vccd1
+ vccd1 _18944_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13018_ _13061_/A vssd1 vssd1 vccd1 vccd1 _13019_/A sky130_fd_sc_hd__buf_2
X_18875_ _19208_/A vssd1 vssd1 vccd1 vccd1 _18875_/X sky130_fd_sc_hd__buf_2
XFILLER_121_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17826_ _18474_/A vssd1 vssd1 vccd1 vccd1 _18379_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17757_ _17757_/A vssd1 vssd1 vccd1 vccd1 _17770_/S sky130_fd_sc_hd__buf_2
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ _15023_/A vssd1 vssd1 vccd1 vccd1 _14981_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16708_ _16708_/A _16708_/B vssd1 vssd1 vccd1 vccd1 _16708_/Y sky130_fd_sc_hd__nand2_1
X_17688_ _17688_/A vssd1 vssd1 vccd1 vccd1 _25915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19427_ _19427_/A vssd1 vssd1 vccd1 vccd1 _26066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16639_ _16639_/A _25907_/Q vssd1 vssd1 vccd1 vccd1 _16640_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19358_ _19492_/A vssd1 vssd1 vccd1 vccd1 _19468_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_176_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18309_ _18398_/A _18309_/B _18309_/C vssd1 vssd1 vccd1 vccd1 _18310_/A sky130_fd_sc_hd__and3_1
XFILLER_200_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19289_ _19286_/X _19288_/X _19334_/S vssd1 vssd1 vccd1 vccd1 _19289_/X sky130_fd_sc_hd__mux2_1
X_21320_ _21320_/A vssd1 vssd1 vccd1 vccd1 _21320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21251_ _21231_/X _21234_/X _21237_/X _21240_/X _21241_/X _21242_/X vssd1 vssd1 vccd1
+ vccd1 _21252_/A sky130_fd_sc_hd__mux4_1
XFILLER_116_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20202_ _20250_/A vssd1 vssd1 vccd1 vccd1 _20202_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21182_ _21214_/A vssd1 vssd1 vccd1 vccd1 _21182_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20133_ _20165_/A vssd1 vssd1 vccd1 vccd1 _20133_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25990_ _26022_/CLK _25990_/D vssd1 vssd1 vccd1 vccd1 _25990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20064_ _20064_/A vssd1 vssd1 vccd1 vccd1 _20064_/X sky130_fd_sc_hd__clkbuf_2
X_24941_ _24941_/A _27777_/Q _24941_/C vssd1 vssd1 vccd1 vccd1 _24947_/B sky130_fd_sc_hd__and3_1
XFILLER_98_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24872_ _27764_/Q _24873_/B vssd1 vssd1 vccd1 vccd1 _24880_/C sky130_fd_sc_hd__and2_1
X_27660_ _27666_/CLK _27660_/D vssd1 vssd1 vccd1 vccd1 _27660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater250 _27604_/CLK vssd1 vssd1 vccd1 vccd1 _27606_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_86_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater261 _27536_/CLK vssd1 vssd1 vccd1 vccd1 _27608_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26611_ _21452_/X _26611_/D vssd1 vssd1 vccd1 vccd1 _26611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23823_ _27072_/Q _23812_/X _23813_/X _27104_/Q _23814_/X vssd1 vssd1 vccd1 vccd1
+ _23823_/X sky130_fd_sc_hd__a221o_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27591_ _27592_/CLK _27591_/D vssd1 vssd1 vccd1 vccd1 _27591_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater272 _27600_/CLK vssd1 vssd1 vccd1 vccd1 _27602_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater283 _27520_/CLK vssd1 vssd1 vccd1 vccd1 _27587_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater294 _27245_/CLK vssd1 vssd1 vccd1 vccd1 _27258_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_306 _24388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26542_ _21206_/X _26542_/D vssd1 vssd1 vccd1 vccd1 _26542_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_317 _24405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23754_ _23777_/A vssd1 vssd1 vccd1 vccd1 _24046_/S sky130_fd_sc_hd__buf_2
XANTENNA_328 _24925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20966_ _20966_/A vssd1 vssd1 vccd1 vccd1 _20966_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_339 _13222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22705_ _22697_/X _22698_/X _22699_/X _22700_/X _22702_/X _22704_/X vssd1 vssd1 vccd1
+ vccd1 _22706_/A sky130_fd_sc_hd__mux4_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26473_ _20968_/X _26473_/D vssd1 vssd1 vccd1 vccd1 _26473_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23685_ _23707_/A vssd1 vssd1 vccd1 vccd1 _23694_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _20886_/X _20888_/X _20890_/X _20892_/X _20893_/X _20894_/X vssd1 vssd1 vccd1
+ vccd1 _20898_/A sky130_fd_sc_hd__mux4_1
XFILLER_0_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25424_ _27750_/Q input62/X _25424_/S vssd1 vssd1 vccd1 vccd1 _25425_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22636_ _22700_/A vssd1 vssd1 vccd1 vccd1 _22636_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25355_ _25355_/A _25355_/B vssd1 vssd1 vccd1 vccd1 _25356_/B sky130_fd_sc_hd__xnor2_1
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22567_ _22561_/X _22562_/X _22563_/X _22564_/X _22565_/X _22566_/X vssd1 vssd1 vccd1
+ vccd1 _22568_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_467 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24306_ _24306_/A _24384_/B vssd1 vssd1 vccd1 vccd1 _27435_/D sky130_fd_sc_hd__nor2_1
X_21518_ _21550_/A vssd1 vssd1 vccd1 vccd1 _21518_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25286_ _27539_/Q _27509_/Q vssd1 vssd1 vccd1 vccd1 _25287_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22498_ _22498_/A vssd1 vssd1 vccd1 vccd1 _22498_/X sky130_fd_sc_hd__clkbuf_1
X_27025_ _22898_/X _27025_/D vssd1 vssd1 vccd1 vccd1 _27025_/Q sky130_fd_sc_hd__dfxtp_1
X_24237_ _24237_/A _24256_/B vssd1 vssd1 vccd1 vccd1 _27390_/D sky130_fd_sc_hd__nor2_1
X_21449_ _21443_/X _21444_/X _21445_/X _21446_/X _21447_/X _21448_/X vssd1 vssd1 vccd1
+ vccd1 _21450_/A sky130_fd_sc_hd__mux4_1
XFILLER_108_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24168_ _24168_/A vssd1 vssd1 vccd1 vccd1 _27355_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23119_ _27101_/Q _17686_/X _23121_/S vssd1 vssd1 vccd1 vccd1 _23120_/A sky130_fd_sc_hd__mux2_1
X_16990_ _27826_/Q _27130_/Q _25875_/Q _25843_/Q _17307_/A _16989_/X vssd1 vssd1 vccd1
+ vccd1 _16990_/X sky130_fd_sc_hd__mux4_1
X_24099_ _24099_/A vssd1 vssd1 vccd1 vccd1 _27324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27927_ _27927_/A _15959_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
X_15941_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15941_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_697 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18660_ _18660_/A vssd1 vssd1 vccd1 vccd1 _25995_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15872_/Y sky130_fd_sc_hd__inv_2
X_27858_ _25808_/X _27858_/D vssd1 vssd1 vccd1 vccd1 _27858_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17611_ _17611_/A vssd1 vssd1 vccd1 vccd1 _25878_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26809_ _22140_/X _26809_/D vssd1 vssd1 vccd1 vccd1 _26809_/Q sky130_fd_sc_hd__dfxtp_1
X_14823_ _14823_/A vssd1 vssd1 vccd1 vccd1 _26518_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _25543_/A vssd1 vssd1 vccd1 vccd1 _18591_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27789_ _27789_/CLK _27789_/D vssd1 vssd1 vccd1 vccd1 _27979_/A sky130_fd_sc_hd__dfxtp_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _17599_/S vssd1 vssd1 vccd1 vccd1 _17551_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14754_ _14753_/X _26540_/Q _14757_/S vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__mux2_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13705_ _13745_/A vssd1 vssd1 vccd1 vccd1 _13705_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17473_ _17505_/A vssd1 vssd1 vccd1 vccd1 _17486_/S sky130_fd_sc_hd__clkbuf_2
X_14685_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14685_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19212_ _19205_/X _19207_/X _19211_/X _19186_/X _19139_/X vssd1 vssd1 vccd1 vccd1
+ _19222_/B sky130_fd_sc_hd__a221o_1
XFILLER_189_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13636_ _13649_/A vssd1 vssd1 vccd1 vccd1 _13647_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_16424_ _16772_/A _16424_/B vssd1 vssd1 vccd1 vccd1 _16479_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19143_ _19261_/A _19143_/B vssd1 vssd1 vccd1 vccd1 _19143_/X sky130_fd_sc_hd__or2_1
XFILLER_81_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13567_ _27338_/Q _13022_/X _13030_/X _27306_/Q _13219_/X vssd1 vssd1 vccd1 vccd1
+ _14521_/A sky130_fd_sc_hd__a221oi_4
X_16355_ _14798_/A _16314_/X _16098_/A _25948_/Q _16354_/Y vssd1 vssd1 vccd1 vccd1
+ _16764_/B sky130_fd_sc_hd__a221o_1
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15306_ _26310_/Q _13382_/X _15306_/S vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16286_ _16801_/A vssd1 vssd1 vccd1 vccd1 _16802_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19074_ _19385_/A vssd1 vssd1 vccd1 vccd1 _19074_/X sky130_fd_sc_hd__clkbuf_2
X_13498_ _13546_/A vssd1 vssd1 vccd1 vccd1 _13517_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18025_ _18023_/X _18024_/X _18075_/S vssd1 vssd1 vccd1 vccd1 _18025_/X sky130_fd_sc_hd__mux2_1
X_15237_ _14775_/X _26341_/Q _15245_/S vssd1 vssd1 vccd1 vccd1 _15238_/A sky130_fd_sc_hd__mux2_1
X_15168_ _15168_/A vssd1 vssd1 vccd1 vccd1 _26372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _26758_/Q _14117_/X _14107_/X _14118_/Y vssd1 vssd1 vccd1 vccd1 _26758_/D
+ sky130_fd_sc_hd__a31o_1
X_15099_ _14785_/X _26402_/Q _15101_/S vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__mux2_1
X_19976_ _19976_/A vssd1 vssd1 vccd1 vccd1 _19976_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18927_ _26141_/Q _26077_/Q _27005_/Q _26973_/Q _18807_/X _24398_/A vssd1 vssd1 vccd1
+ vccd1 _18928_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ _19004_/A _18858_/B vssd1 vssd1 vccd1 vccd1 _18858_/X sky130_fd_sc_hd__or2_1
XFILLER_80_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17809_ _27594_/Q vssd1 vssd1 vccd1 vccd1 _18182_/A sky130_fd_sc_hd__clkbuf_2
X_18789_ _19460_/A vssd1 vssd1 vccd1 vccd1 _19412_/A sky130_fd_sc_hd__buf_2
X_20820_ _20852_/A vssd1 vssd1 vccd1 vccd1 _20820_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20751_ _20751_/A vssd1 vssd1 vccd1 vccd1 _20751_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23470_ _27181_/Q _23470_/B vssd1 vssd1 vccd1 vccd1 _23470_/X sky130_fd_sc_hd__or2_1
XFILLER_196_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20682_ _20668_/X _20669_/X _20670_/X _20671_/X _20672_/X _20673_/X vssd1 vssd1 vccd1
+ vccd1 _20683_/A sky130_fd_sc_hd__mux4_1
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22421_ _22421_/A vssd1 vssd1 vccd1 vccd1 _22421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25140_ _27693_/Q _25112_/X _25139_/Y _25132_/X vssd1 vssd1 vccd1 vccd1 _27693_/D
+ sky130_fd_sc_hd__o211a_1
X_22352_ _22421_/A vssd1 vssd1 vccd1 vccd1 _22352_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21303_ _21303_/A vssd1 vssd1 vccd1 vccd1 _21303_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25071_ _25923_/Q _25989_/Q _25822_/Q _26021_/Q _25052_/X _25070_/X vssd1 vssd1 vccd1
+ vccd1 _25071_/X sky130_fd_sc_hd__mux4_1
X_22283_ _22455_/A vssd1 vssd1 vccd1 vccd1 _22349_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24022_ _27854_/Q _27158_/Q _25903_/Q _25871_/Q _24014_/X _23991_/X vssd1 vssd1 vccd1
+ vccd1 _24022_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21234_ _21302_/A vssd1 vssd1 vccd1 vccd1 _21234_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21165_ _21213_/A vssd1 vssd1 vccd1 vccd1 _21165_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20116_ _20164_/A vssd1 vssd1 vccd1 vccd1 _20116_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25973_ _25974_/CLK _25973_/D vssd1 vssd1 vccd1 vccd1 _25973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21096_ _21128_/A vssd1 vssd1 vccd1 vccd1 _21096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27712_ _27770_/CLK _27712_/D vssd1 vssd1 vccd1 vccd1 _27712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20047_ _20079_/A vssd1 vssd1 vccd1 vccd1 _20047_/X sky130_fd_sc_hd__clkbuf_1
X_24924_ _27661_/Q _24909_/X _24923_/Y _24914_/X vssd1 vssd1 vccd1 vccd1 _27661_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27643_ _27753_/CLK _27643_/D vssd1 vssd1 vccd1 vccd1 _27643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24855_ _27647_/Q _24834_/X _24854_/Y _24839_/X vssd1 vssd1 vccd1 vccd1 _27647_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_435 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _19419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_114 _22537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23806_ _24045_/S vssd1 vssd1 vccd1 vccd1 _23844_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _22616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24786_ _24786_/A _24786_/B vssd1 vssd1 vccd1 vccd1 _24786_/Y sky130_fd_sc_hd__nand2_1
X_27574_ _27574_/CLK _27574_/D vssd1 vssd1 vccd1 vccd1 _27574_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _21998_/A vssd1 vssd1 vccd1 vccd1 _21998_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _23598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _13105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26525_ _21154_/X _26525_/D vssd1 vssd1 vccd1 vccd1 _26525_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_158 _13379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23737_ _23737_/A vssd1 vssd1 vccd1 vccd1 _27270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20949_ _20937_/X _20938_/X _20939_/X _20940_/X _20941_/X _20942_/X vssd1 vssd1 vccd1
+ vccd1 _20950_/A sky130_fd_sc_hd__mux4_1
XFILLER_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_169 _13414_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14470_ _26636_/Q _14460_/X _14455_/X _14469_/Y vssd1 vssd1 vccd1 vccd1 _26636_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26456_ _20914_/X _26456_/D vssd1 vssd1 vccd1 vccd1 _26456_/Q sky130_fd_sc_hd__dfxtp_1
X_23668_ _27760_/Q _27240_/Q _23672_/S vssd1 vssd1 vccd1 vccd1 _23669_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ _26970_/Q _13420_/X _13421_/S vssd1 vssd1 vccd1 vccd1 _13422_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22619_ _22609_/X _22610_/X _22611_/X _22612_/X _22615_/X _22618_/X vssd1 vssd1 vccd1
+ vccd1 _22620_/A sky130_fd_sc_hd__mux4_1
X_25407_ _27742_/Q input54/X _25413_/S vssd1 vssd1 vccd1 vccd1 _25408_/A sky130_fd_sc_hd__mux2_1
X_26387_ _20663_/X _26387_/D vssd1 vssd1 vccd1 vccd1 _26387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23599_ _27778_/Q vssd1 vssd1 vccd1 vccd1 _24941_/A sky130_fd_sc_hd__buf_2
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16140_ _26069_/Q _16137_/X _16139_/X vssd1 vssd1 vccd1 vccd1 _24306_/A sky130_fd_sc_hd__a21oi_2
X_25338_ _25347_/A _27515_/Q vssd1 vssd1 vccd1 vccd1 _25339_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _13352_/A vssd1 vssd1 vccd1 vccd1 _26992_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16071_ _27407_/Q _16094_/A vssd1 vssd1 vccd1 vccd1 _16071_/Y sky130_fd_sc_hd__nand2_1
X_25269_ _27539_/Q vssd1 vssd1 vccd1 vccd1 _25323_/A sky130_fd_sc_hd__clkbuf_4
X_13283_ _27018_/Q _13144_/X _13291_/S vssd1 vssd1 vccd1 vccd1 _13284_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15022_ _26435_/Q _15015_/X _15016_/X _15021_/Y vssd1 vssd1 vccd1 vccd1 _26435_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27008_ _22834_/X _27008_/D vssd1 vssd1 vccd1 vccd1 _27008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19830_ _19830_/A vssd1 vssd1 vccd1 vccd1 _19898_/A sky130_fd_sc_hd__buf_2
XFILLER_150_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19761_ _19761_/A vssd1 vssd1 vccd1 vccd1 _19761_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16973_ _16973_/A vssd1 vssd1 vccd1 vccd1 _25911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18712_ _18712_/A vssd1 vssd1 vccd1 vccd1 _26018_/D sky130_fd_sc_hd__clkbuf_1
X_15924_ _15924_/A vssd1 vssd1 vccd1 vccd1 _15924_/Y sky130_fd_sc_hd__inv_2
X_19692_ _19678_/X _19679_/X _19680_/X _19681_/X _19682_/X _19683_/X vssd1 vssd1 vccd1
+ vccd1 _19693_/A sky130_fd_sc_hd__mux4_1
Xinput9 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_188_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18643_ _18689_/S vssd1 vssd1 vccd1 vccd1 _18652_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ input1/X vssd1 vssd1 vccd1 vccd1 _15980_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _14806_/A vssd1 vssd1 vccd1 vccd1 _26524_/D sky130_fd_sc_hd__clkbuf_1
X_18574_ _26169_/Q _26105_/Q _27033_/Q _27001_/Q _17810_/X _18011_/X vssd1 vssd1 vccd1
+ vccd1 _18575_/A sky130_fd_sc_hd__mux4_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15786_ _13038_/X _26105_/Q _15794_/S vssd1 vssd1 vccd1 vccd1 _15787_/A sky130_fd_sc_hd__mux2_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12998_ _27799_/Q _12998_/B vssd1 vssd1 vccd1 vccd1 _12999_/A sky130_fd_sc_hd__and2_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17525_ _17525_/A vssd1 vssd1 vccd1 vccd1 _25842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14737_ _14737_/A vssd1 vssd1 vccd1 vccd1 _14737_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17456_ _27418_/Q vssd1 vssd1 vccd1 vccd1 _17456_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14668_ _26570_/Q _14658_/X _14666_/X _14667_/Y vssd1 vssd1 vccd1 vccd1 _26570_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ _16407_/A vssd1 vssd1 vccd1 vccd1 _16447_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13619_ _13889_/A _13621_/B vssd1 vssd1 vccd1 vccd1 _13619_/Y sky130_fd_sc_hd__nor2_1
X_17387_ _27226_/Q _17386_/X _17387_/S vssd1 vssd1 vccd1 vccd1 _17388_/A sky130_fd_sc_hd__mux2_1
X_14599_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14610_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19126_ _26405_/Q _26373_/Q _26341_/Q _26309_/Q _19054_/X _19100_/X vssd1 vssd1 vccd1
+ vccd1 _19126_/X sky130_fd_sc_hd__mux4_1
XFILLER_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16338_ _16266_/A _16182_/X _16185_/X _16186_/X vssd1 vssd1 vccd1 vccd1 _16759_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19057_ _19055_/X _19056_/X _19057_/S vssd1 vssd1 vccd1 vccd1 _19057_/X sky130_fd_sc_hd__mux2_1
X_16269_ _27393_/Q vssd1 vssd1 vccd1 vccd1 _16490_/A sky130_fd_sc_hd__inv_2
XFILLER_69_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18008_ _18008_/A _24392_/A vssd1 vssd1 vccd1 vccd1 _18008_/X sky130_fd_sc_hd__or2b_1
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19959_ _19991_/A vssd1 vssd1 vccd1 vccd1 _19959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28013__479 vssd1 vssd1 vccd1 vccd1 _28013__479/HI _28013_/A sky130_fd_sc_hd__conb_1
X_22970_ _22970_/A vssd1 vssd1 vccd1 vccd1 _22970_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21921_ _21911_/X _21912_/X _21913_/X _21914_/X _21916_/X _21918_/X vssd1 vssd1 vccd1
+ vccd1 _21922_/A sky130_fd_sc_hd__mux4_1
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24640_ _24640_/A _25110_/B vssd1 vssd1 vccd1 vccd1 _24748_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21852_ _21900_/A vssd1 vssd1 vccd1 vccd1 _21852_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20803_ _20867_/A vssd1 vssd1 vccd1 vccd1 _20803_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24571_ _24571_/A vssd1 vssd1 vccd1 vccd1 _27546_/D sky130_fd_sc_hd__clkbuf_1
X_21783_ _21777_/X _21778_/X _21779_/X _21780_/X _21781_/X _21782_/X vssd1 vssd1 vccd1
+ vccd1 _21784_/A sky130_fd_sc_hd__mux4_1
XFILLER_24_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26310_ _20399_/X _26310_/D vssd1 vssd1 vccd1 vccd1 _26310_/Q sky130_fd_sc_hd__dfxtp_1
X_23522_ _23526_/A _23522_/B vssd1 vssd1 vccd1 vccd1 _23523_/A sky130_fd_sc_hd__and2_1
X_27290_ _27786_/CLK _27290_/D vssd1 vssd1 vccd1 vccd1 _27290_/Q sky130_fd_sc_hd__dfxtp_1
X_20734_ _20722_/X _20723_/X _20724_/X _20725_/X _20726_/X _20727_/X vssd1 vssd1 vccd1
+ vccd1 _20735_/A sky130_fd_sc_hd__mux4_1
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26241_ _20155_/X _26241_/D vssd1 vssd1 vccd1 vccd1 _26241_/Q sky130_fd_sc_hd__dfxtp_1
X_23453_ _27175_/Q _23456_/B vssd1 vssd1 vccd1 vccd1 _23453_/X sky130_fd_sc_hd__or2_1
XFILLER_17_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20665_ _20665_/A vssd1 vssd1 vccd1 vccd1 _20665_/X sky130_fd_sc_hd__clkbuf_1
X_22404_ _22436_/A vssd1 vssd1 vccd1 vccd1 _22404_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26172_ _19911_/X _26172_/D vssd1 vssd1 vccd1 vccd1 _26172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23384_ _27776_/Q vssd1 vssd1 vccd1 vccd1 _24794_/A sky130_fd_sc_hd__inv_2
XFILLER_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20596_ _20582_/X _20583_/X _20584_/X _20585_/X _20586_/X _20587_/X vssd1 vssd1 vccd1
+ vccd1 _20597_/A sky130_fd_sc_hd__mux4_2
XFILLER_137_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25123_ _25139_/A _25123_/B vssd1 vssd1 vccd1 vccd1 _25123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22335_ _22335_/A vssd1 vssd1 vccd1 vccd1 _22335_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25054_ _27231_/Q vssd1 vssd1 vccd1 vccd1 _25087_/S sky130_fd_sc_hd__clkbuf_2
X_22266_ _22335_/A vssd1 vssd1 vccd1 vccd1 _22266_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24005_ _24005_/A vssd1 vssd1 vccd1 vccd1 _24005_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21217_ _21217_/A vssd1 vssd1 vccd1 vccd1 _21290_/A sky130_fd_sc_hd__clkbuf_2
X_22197_ _22455_/A vssd1 vssd1 vccd1 vccd1 _22263_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21148_ _21213_/A vssd1 vssd1 vccd1 vccd1 _21148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13970_ _16298_/A vssd1 vssd1 vccd1 vccd1 _14348_/A sky130_fd_sc_hd__buf_2
XFILLER_120_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21079_ _21127_/A vssd1 vssd1 vccd1 vccd1 _21079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25956_ _26057_/CLK _25956_/D vssd1 vssd1 vccd1 vccd1 _25956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _12921_/A _12921_/B vssd1 vssd1 vccd1 vccd1 _12929_/A sky130_fd_sc_hd__nand2_1
X_24907_ _24913_/A _24907_/B vssd1 vssd1 vccd1 vccd1 _24907_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25887_ _27141_/CLK _25887_/D vssd1 vssd1 vccd1 vccd1 _25887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27626_ _27627_/CLK _27626_/D vssd1 vssd1 vccd1 vccd1 _27626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15640_ _15640_/A vssd1 vssd1 vccd1 vccd1 _26163_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24838_ _24838_/A _24838_/B vssd1 vssd1 vccd1 vccd1 _24838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27557_ _27558_/CLK _27557_/D vssd1 vssd1 vccd1 vccd1 _27557_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _26193_/Q _14737_/A _15573_/S vssd1 vssd1 vccd1 vccd1 _15572_/A sky130_fd_sc_hd__mux2_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24769_ _24769_/A _24772_/B vssd1 vssd1 vccd1 vccd1 _24769_/Y sky130_fd_sc_hd__nand2_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17306_/X _17308_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17310_/X sky130_fd_sc_hd__mux2_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _15775_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14522_/Y sky130_fd_sc_hd__nor2_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26508_ _21090_/X _26508_/D vssd1 vssd1 vccd1 vccd1 _26508_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18290_ _26956_/Q _26924_/Q _26892_/Q _26860_/Q _17999_/X _18000_/X vssd1 vssd1 vccd1
+ vccd1 _18290_/X sky130_fd_sc_hd__mux4_2
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27488_ _27488_/CLK _27488_/D vssd1 vssd1 vccd1 vccd1 _27488_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17216_/X _17241_/B vssd1 vssd1 vccd1 vccd1 _17241_/X sky130_fd_sc_hd__and2b_1
XFILLER_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14453_ _15725_/A _14465_/B vssd1 vssd1 vccd1 vccd1 _14453_/Y sky130_fd_sc_hd__nor2_1
X_26439_ _20847_/X _26439_/D vssd1 vssd1 vccd1 vccd1 _26439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13404_ _13404_/A vssd1 vssd1 vccd1 vccd1 _26976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14384_ _26662_/Q _14379_/X _14371_/X _14383_/Y vssd1 vssd1 vccd1 vccd1 _26662_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_167_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17172_ _17116_/X _17166_/X _17168_/X _17171_/X vssd1 vssd1 vccd1 vccd1 _17172_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_167_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16123_ _16111_/Y _16119_/X _16121_/X _16099_/A _16122_/Y vssd1 vssd1 vccd1 vccd1
+ _24309_/A sky130_fd_sc_hd__o221a_2
X_13335_ _26997_/Q _13334_/X _13335_/S vssd1 vssd1 vccd1 vccd1 _13336_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16054_ _16052_/Y _16017_/B _16014_/B _16053_/Y vssd1 vssd1 vccd1 vccd1 _16054_/X
+ sky130_fd_sc_hd__a22o_1
X_13266_ _13266_/A vssd1 vssd1 vccd1 vccd1 _27026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15005_ _26442_/Q _15002_/X _15003_/X _15004_/Y vssd1 vssd1 vccd1 vccd1 _26442_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13197_ _27342_/Q _13193_/X _13194_/X _27310_/Q _13196_/X vssd1 vssd1 vccd1 vccd1
+ _16206_/A sky130_fd_sc_hd__a221o_4
XFILLER_123_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19813_ _19813_/A vssd1 vssd1 vccd1 vccd1 _19813_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19744_ _19830_/A vssd1 vssd1 vccd1 vccd1 _19812_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16956_ _24635_/B _24626_/D vssd1 vssd1 vccd1 vccd1 _24488_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15907_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15912_/A sky130_fd_sc_hd__buf_2
XFILLER_65_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_593 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19675_ _19675_/A vssd1 vssd1 vccd1 vccd1 _19675_/X sky130_fd_sc_hd__clkbuf_1
X_16887_ _16077_/A _16798_/A _16798_/B _16621_/X vssd1 vssd1 vccd1 vccd1 _16887_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_2_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18626_ _25980_/Q _17683_/X _18630_/S vssd1 vssd1 vccd1 vccd1 _18627_/A sky130_fd_sc_hd__mux2_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _13198_/X _26081_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15839_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18557_ _18557_/A _18479_/X vssd1 vssd1 vccd1 vccd1 _18557_/X sky130_fd_sc_hd__or2b_1
X_15769_ _15769_/A _15771_/B vssd1 vssd1 vccd1 vccd1 _15769_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17508_ _27434_/Q vssd1 vssd1 vccd1 vccd1 _17508_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18488_ _18485_/X _18487_/X _18488_/S vssd1 vssd1 vccd1 vccd1 _18488_/X sky130_fd_sc_hd__mux2_2
XFILLER_162_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_14 _25926_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17439_ _17439_/A vssd1 vssd1 vccd1 vccd1 _25815_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_25 _27141_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 _18458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _17970_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 _18245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20450_ _20708_/A vssd1 vssd1 vccd1 vccd1 _20515_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_69 _18344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19109_ _19473_/A vssd1 vssd1 vccd1 vccd1 _19222_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20381_ _20413_/A vssd1 vssd1 vccd1 vccd1 _20381_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22120_ _22120_/A vssd1 vssd1 vccd1 vccd1 _22120_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22051_ _22083_/A vssd1 vssd1 vccd1 vccd1 _22051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21002_ _21002_/A vssd1 vssd1 vccd1 vccd1 _21002_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25810_ _25810_/A vssd1 vssd1 vccd1 vccd1 _25810_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26790_ _22074_/X _26790_/D vssd1 vssd1 vccd1 vccd1 _26790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22953_ _22939_/X _22940_/X _22941_/X _22942_/X _22943_/X _22944_/X vssd1 vssd1 vccd1
+ vccd1 _22954_/A sky130_fd_sc_hd__mux4_1
X_25741_ _25741_/A vssd1 vssd1 vccd1 vccd1 _27827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21904_ _21904_/A vssd1 vssd1 vccd1 vccd1 _21904_/X sky130_fd_sc_hd__clkbuf_1
X_25672_ _25672_/A vssd1 vssd1 vccd1 vccd1 _25672_/X sky130_fd_sc_hd__clkbuf_1
X_22884_ _22884_/A vssd1 vssd1 vccd1 vccd1 _22884_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27411_ _27411_/CLK _27411_/D vssd1 vssd1 vccd1 vccd1 _27411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21835_ _21825_/X _21826_/X _21827_/X _21828_/X _21830_/X _21832_/X vssd1 vssd1 vccd1
+ vccd1 _21836_/A sky130_fd_sc_hd__mux4_1
X_24623_ _24623_/A vssd1 vssd1 vccd1 vccd1 _27570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24554_ _24554_/A _24554_/B vssd1 vssd1 vccd1 vccd1 _24555_/A sky130_fd_sc_hd__and2_1
X_27342_ _27342_/CLK _27342_/D vssd1 vssd1 vccd1 vccd1 _27342_/Q sky130_fd_sc_hd__dfxtp_2
X_21766_ _21814_/A vssd1 vssd1 vccd1 vccd1 _21766_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20717_ _20717_/A vssd1 vssd1 vccd1 vccd1 _20717_/X sky130_fd_sc_hd__clkbuf_1
X_23505_ _23415_/X _23503_/X _25430_/B vssd1 vssd1 vccd1 vccd1 _27194_/D sky130_fd_sc_hd__a21o_1
X_24485_ _27639_/Q _24509_/B vssd1 vssd1 vccd1 vccd1 _24486_/A sky130_fd_sc_hd__and2_1
X_27273_ _27379_/CLK _27273_/D vssd1 vssd1 vccd1 vccd1 _27273_/Q sky130_fd_sc_hd__dfxtp_1
X_21697_ _21689_/X _21690_/X _21691_/X _21692_/X _21693_/X _21694_/X vssd1 vssd1 vccd1
+ vccd1 _21698_/A sky130_fd_sc_hd__mux4_1
XFILLER_200_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23436_ _27168_/Q _23443_/B vssd1 vssd1 vccd1 vccd1 _23436_/X sky130_fd_sc_hd__or2_1
X_26224_ _20093_/X _26224_/D vssd1 vssd1 vccd1 vccd1 _26224_/Q sky130_fd_sc_hd__dfxtp_1
X_20648_ _20636_/X _20637_/X _20638_/X _20639_/X _20640_/X _20641_/X vssd1 vssd1 vccd1
+ vccd1 _20649_/A sky130_fd_sc_hd__mux4_1
XFILLER_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26155_ _19857_/X _26155_/D vssd1 vssd1 vccd1 vccd1 _26155_/Q sky130_fd_sc_hd__dfxtp_1
X_23367_ _24792_/A _27255_/Q _27248_/Q _24772_/A vssd1 vssd1 vccd1 vccd1 _23367_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_20579_ _20579_/A vssd1 vssd1 vccd1 vccd1 _20579_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13120_ _27291_/Q _13125_/B vssd1 vssd1 vccd1 vccd1 _13120_/X sky130_fd_sc_hd__and2_2
X_22318_ _22350_/A vssd1 vssd1 vccd1 vccd1 _22318_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25106_ _25106_/A _25110_/B vssd1 vssd1 vccd1 vccd1 _25107_/A sky130_fd_sc_hd__and2_1
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26086_ _19614_/X _26086_/D vssd1 vssd1 vccd1 vccd1 _26086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23298_ _23272_/Y input44/X _27736_/Q _23295_/Y _23297_/X vssd1 vssd1 vccd1 vccd1
+ _23300_/B sky130_fd_sc_hd__a221o_1
XFILLER_30_1182 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _13241_/S vssd1 vssd1 vccd1 vccd1 _13079_/S sky130_fd_sc_hd__clkbuf_2
X_25037_ _25919_/Q _25985_/Q _25818_/Q _26017_/Q _25009_/X _25027_/X vssd1 vssd1 vccd1
+ vccd1 _25037_/X sky130_fd_sc_hd__mux4_1
X_22249_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22249_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16810_ _16666_/Y _16665_/X _16809_/Y vssd1 vssd1 vccd1 vccd1 _16811_/D sky130_fd_sc_hd__o21a_1
XFILLER_120_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17790_ _18455_/A vssd1 vssd1 vccd1 vccd1 _18425_/A sky130_fd_sc_hd__buf_2
XFILLER_8_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26988_ _22764_/X _26988_/D vssd1 vssd1 vccd1 vccd1 _26988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16741_ _16737_/X _16738_/Y _16740_/Y vssd1 vssd1 vccd1 vccd1 _24225_/A sky130_fd_sc_hd__o21a_1
XFILLER_98_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25939_ _27855_/CLK _25939_/D vssd1 vssd1 vccd1 vccd1 _25939_/Q sky130_fd_sc_hd__dfxtp_1
X_13953_ _14425_/A vssd1 vssd1 vccd1 vccd1 _14335_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19460_ _19460_/A vssd1 vssd1 vccd1 vccd1 _19460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672_ _16672_/A _16672_/B vssd1 vssd1 vccd1 vccd1 _16672_/Y sky130_fd_sc_hd__xnor2_1
X_13884_ _13884_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13884_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _18379_/X _18407_/X _18410_/X _18384_/X vssd1 vssd1 vccd1 vccd1 _18411_/X
+ sky130_fd_sc_hd__o211a_1
X_27609_ _27611_/CLK _27609_/D vssd1 vssd1 vccd1 vccd1 _27609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15623_ _15783_/A _15623_/B vssd1 vssd1 vccd1 vccd1 _15680_/A sky130_fd_sc_hd__or2_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _19391_/A vssd1 vssd1 vccd1 vccd1 _19480_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18336_/X _18338_/X _18341_/X _18468_/A vssd1 vssd1 vccd1 vccd1 _18342_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _26201_/Q _14709_/A _15562_/S vssd1 vssd1 vccd1 vccd1 _15555_/A sky130_fd_sc_hd__mux2_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _15762_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14505_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _26699_/Q _26667_/Q _26635_/Q _26603_/Q _18177_/X _18249_/X vssd1 vssd1 vccd1
+ vccd1 _18274_/A sky130_fd_sc_hd__mux4_1
XFILLER_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15485_ _15485_/A vssd1 vssd1 vccd1 vccd1 _26232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17224_ _17222_/X _17223_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17224_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14436_ _14436_/A vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 la1_data_in[12] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_6
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 la1_data_in[22] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_4
XFILLER_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 la1_data_in[3] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17155_ _17338_/A vssd1 vssd1 vccd1 vccd1 _17155_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput45 la1_oenb[13] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_8
X_14367_ _14367_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14367_/Y sky130_fd_sc_hd__nor2_1
Xinput56 la1_oenb[23] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_6
XFILLER_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput67 la1_oenb[4] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_4
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16106_ _16106_/A vssd1 vssd1 vccd1 vccd1 _16576_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13318_ _13318_/A vssd1 vssd1 vccd1 vccd1 _27002_/D sky130_fd_sc_hd__clkbuf_1
X_14298_ _14386_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14298_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17086_ _25817_/Q _26016_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17086_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16037_ _16026_/X _16029_/Y _16033_/X _16036_/X vssd1 vssd1 vccd1 vccd1 _16845_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13249_ _13317_/S vssd1 vssd1 vccd1 vccd1 _13258_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17988_ _26399_/Q _26367_/Q _26335_/Q _26303_/Q _17877_/X _17943_/X vssd1 vssd1 vccd1
+ vccd1 _17988_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19727_ _19727_/A vssd1 vssd1 vccd1 vccd1 _19727_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16939_ _27602_/Q _27488_/Q vssd1 vssd1 vccd1 vccd1 _16945_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19658_ _19830_/A vssd1 vssd1 vccd1 vccd1 _19726_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18609_ _18589_/X _18600_/X _18604_/Y _18608_/Y vssd1 vssd1 vccd1 vccd1 _25976_/D
+ sky130_fd_sc_hd__o211a_1
X_19589_ _19637_/A vssd1 vssd1 vccd1 vccd1 _19589_/X sky130_fd_sc_hd__clkbuf_1
X_21620_ _21636_/A vssd1 vssd1 vccd1 vccd1 _21620_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21551_ _21545_/X _21546_/X _21547_/X _21548_/X _21549_/X _21550_/X vssd1 vssd1 vccd1
+ vccd1 _21552_/A sky130_fd_sc_hd__mux4_1
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20502_ _20496_/X _20497_/X _20498_/X _20499_/X _20500_/X _20501_/X vssd1 vssd1 vccd1
+ vccd1 _20503_/A sky130_fd_sc_hd__mux4_1
X_24270_ _16182_/X _16185_/X _24269_/X vssd1 vssd1 vccd1 vccd1 _27408_/D sky130_fd_sc_hd__o21a_1
X_21482_ _21550_/A vssd1 vssd1 vccd1 vccd1 _21482_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23221_ _23221_/A vssd1 vssd1 vccd1 vccd1 _27146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20433_ _20501_/A vssd1 vssd1 vccd1 vccd1 _20433_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23152_ _27116_/Q _17734_/X _23154_/S vssd1 vssd1 vccd1 vccd1 _23153_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20364_ _20412_/A vssd1 vssd1 vccd1 vccd1 _20364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22103_ _22173_/A vssd1 vssd1 vccd1 vccd1 _22103_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23083_ _23094_/A vssd1 vssd1 vccd1 vccd1 _23092_/S sky130_fd_sc_hd__clkbuf_2
X_27960_ _27960_/A _15871_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20295_ _20295_/A vssd1 vssd1 vccd1 vccd1 _20295_/X sky130_fd_sc_hd__clkbuf_1
X_28019__485 vssd1 vssd1 vccd1 vccd1 _28019__485/HI _28019_/A sky130_fd_sc_hd__conb_1
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22034_ _22034_/A vssd1 vssd1 vccd1 vccd1 _22034_/X sky130_fd_sc_hd__clkbuf_1
X_26911_ _22496_/X _26911_/D vssd1 vssd1 vccd1 vccd1 _26911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26842_ _22256_/X _26842_/D vssd1 vssd1 vccd1 vccd1 _26842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26773_ _22012_/X _26773_/D vssd1 vssd1 vccd1 vccd1 _26773_/Q sky130_fd_sc_hd__dfxtp_1
X_23985_ _23983_/X _23984_/X _23985_/S vssd1 vssd1 vccd1 vccd1 _23985_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25724_ _25724_/A vssd1 vssd1 vccd1 vccd1 _25724_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22936_ _22936_/A vssd1 vssd1 vccd1 vccd1 _22936_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25655_ _25655_/A vssd1 vssd1 vccd1 vccd1 _25722_/A sky130_fd_sc_hd__clkbuf_2
X_22867_ _22853_/X _22854_/X _22855_/X _22856_/X _22857_/X _22858_/X vssd1 vssd1 vccd1
+ vccd1 _22868_/A sky130_fd_sc_hd__mux4_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24606_ _24606_/A vssd1 vssd1 vccd1 vccd1 _27562_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21818_ _21818_/A vssd1 vssd1 vccd1 vccd1 _21818_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25586_ _25560_/X _25313_/B _25585_/X _25566_/X vssd1 vssd1 vccd1 vccd1 _25586_/X
+ sky130_fd_sc_hd__a211o_1
X_22798_ _22798_/A vssd1 vssd1 vccd1 vccd1 _22798_/X sky130_fd_sc_hd__clkbuf_1
X_27325_ _27325_/CLK _27325_/D vssd1 vssd1 vccd1 vccd1 _27325_/Q sky130_fd_sc_hd__dfxtp_1
X_21749_ _21737_/X _21738_/X _21739_/X _21740_/X _21743_/X _21746_/X vssd1 vssd1 vccd1
+ vccd1 _21750_/A sky130_fd_sc_hd__mux4_1
X_24537_ _24537_/A vssd1 vssd1 vccd1 vccd1 _27533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27256_ _27782_/CLK _27256_/D vssd1 vssd1 vccd1 vccd1 _27256_/Q sky130_fd_sc_hd__dfxtp_1
X_15270_ _15270_/A vssd1 vssd1 vccd1 vccd1 _26327_/D sky130_fd_sc_hd__clkbuf_1
X_24468_ _24468_/A vssd1 vssd1 vccd1 vccd1 _27510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14221_ _14399_/A _14226_/B vssd1 vssd1 vccd1 vccd1 _14221_/Y sky130_fd_sc_hd__nor2_1
X_26207_ _20039_/X _26207_/D vssd1 vssd1 vccd1 vccd1 _26207_/Q sky130_fd_sc_hd__dfxtp_1
X_23419_ _27162_/Q _23430_/B vssd1 vssd1 vccd1 vccd1 _23419_/X sky130_fd_sc_hd__or2_1
X_27187_ _27729_/CLK _27187_/D vssd1 vssd1 vccd1 vccd1 _27187_/Q sky130_fd_sc_hd__dfxtp_1
X_24399_ _24399_/A vssd1 vssd1 vccd1 vccd1 _27479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _14166_/A vssd1 vssd1 vccd1 vccd1 _14158_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26138_ _19793_/X _26138_/D vssd1 vssd1 vccd1 vccd1 _26138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13103_ _27294_/Q _13125_/B vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__and2_2
XFILLER_113_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14083_ _14348_/A _14085_/B vssd1 vssd1 vccd1 vccd1 _14083_/Y sky130_fd_sc_hd__nor2_1
X_18960_ _26398_/Q _26366_/Q _26334_/Q _26302_/Q _18887_/X _18826_/X vssd1 vssd1 vccd1
+ vccd1 _18960_/X sky130_fd_sc_hd__mux4_1
X_26069_ _26069_/CLK _26069_/D vssd1 vssd1 vccd1 vccd1 _26069_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _13176_/B vssd1 vssd1 vccd1 vccd1 _13169_/B sky130_fd_sc_hd__clkbuf_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _17911_/A _17910_/X vssd1 vssd1 vccd1 vccd1 _17911_/X sky130_fd_sc_hd__or2b_1
XFILLER_191_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18891_ _18884_/X _18886_/X _18890_/X _18866_/X _18840_/X vssd1 vssd1 vccd1 vccd1
+ _18892_/C sky130_fd_sc_hd__a221o_1
XFILLER_6_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17842_ _17900_/A vssd1 vssd1 vccd1 vccd1 _18141_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17773_ _25942_/Q _17772_/X _17776_/S vssd1 vssd1 vccd1 vccd1 _17774_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14985_ _26449_/Q _14974_/X _14976_/X _14984_/Y vssd1 vssd1 vccd1 vccd1 _26449_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19512_ _19506_/X _19508_/X _19511_/X _19448_/X _19469_/X vssd1 vssd1 vccd1 vccd1
+ _19513_/C sky130_fd_sc_hd__a221o_1
X_16724_ _16619_/A _16890_/C _16719_/Y _16723_/X vssd1 vssd1 vccd1 vccd1 _24231_/A
+ sky130_fd_sc_hd__a31oi_1
X_13936_ _13936_/A _13940_/B vssd1 vssd1 vccd1 vccd1 _13936_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19443_ _19351_/X _19442_/X _19354_/X vssd1 vssd1 vccd1 vccd1 _19443_/X sky130_fd_sc_hd__o21a_1
X_16655_ _16647_/X _16648_/X _16650_/Y _16654_/Y _16877_/A vssd1 vssd1 vccd1 vccd1
+ _24258_/A sky130_fd_sc_hd__o32a_1
XFILLER_62_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13867_ _13920_/A vssd1 vssd1 vccd1 vccd1 _13878_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15606_ _26177_/Q _16206_/A _15606_/S vssd1 vssd1 vccd1 vccd1 _15607_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19374_ _26544_/Q _26512_/Q _26480_/Q _27056_/Q _18926_/A _18923_/X vssd1 vssd1 vccd1
+ vccd1 _19374_/X sky130_fd_sc_hd__mux4_1
X_16586_ _16578_/Y _16584_/Y _16913_/B vssd1 vssd1 vccd1 vccd1 _16586_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _26862_/Q _13793_/X _13794_/X _13797_/Y vssd1 vssd1 vccd1 vccd1 _26862_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_163_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18325_ _26285_/Q _26253_/Q _26221_/Q _26189_/Q _18301_/X _18324_/X vssd1 vssd1 vccd1
+ vccd1 _18325_/X sky130_fd_sc_hd__mux4_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15537_ _13204_/X _26208_/Q _15545_/S vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18256_ _18256_/A _18207_/X vssd1 vssd1 vccd1 vccd1 _18256_/X sky130_fd_sc_hd__or2b_1
XFILLER_176_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15468_ _15468_/A vssd1 vssd1 vccd1 vccd1 _26239_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17207_ _17155_/X _17207_/B vssd1 vssd1 vccd1 vccd1 _17207_/X sky130_fd_sc_hd__and2b_1
X_14419_ _15699_/A _14426_/B vssd1 vssd1 vccd1 vccd1 _14419_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18187_ _18162_/X _18186_/X _18070_/X vssd1 vssd1 vccd1 vccd1 _18187_/X sky130_fd_sc_hd__o21a_1
XFILLER_190_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15399_ _14801_/X _26269_/Q _15401_/S vssd1 vssd1 vccd1 vccd1 _15400_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17138_ _17136_/X _17137_/X _17174_/S vssd1 vssd1 vccd1 vccd1 _17138_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17069_ _17252_/A vssd1 vssd1 vccd1 vccd1 _17069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20080_ _20338_/A vssd1 vssd1 vccd1 vccd1 _20150_/A sky130_fd_sc_hd__buf_2
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater410 _26051_/CLK vssd1 vssd1 vccd1 vccd1 _26048_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater421 _27323_/CLK vssd1 vssd1 vccd1 vccd1 _27331_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater432 _17407_/Y vssd1 vssd1 vccd1 vccd1 _25963_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23770_ _27827_/Q _27131_/Q _25876_/Q _25844_/Q _23997_/A _23744_/X vssd1 vssd1 vccd1
+ vccd1 _23770_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20982_ _20982_/A vssd1 vssd1 vccd1 vccd1 _20982_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22721_ _22893_/A vssd1 vssd1 vccd1 vccd1 _22786_/A sky130_fd_sc_hd__buf_2
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22652_ _22700_/A vssd1 vssd1 vccd1 vccd1 _22652_/X sky130_fd_sc_hd__clkbuf_1
X_25440_ _25552_/A vssd1 vssd1 vccd1 vccd1 _25440_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21603_ _21635_/A vssd1 vssd1 vccd1 vccd1 _21603_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22583_ _22577_/X _22578_/X _22579_/X _22580_/X _22581_/X _22582_/X vssd1 vssd1 vccd1
+ vccd1 _22584_/A sky130_fd_sc_hd__mux4_1
X_25371_ _25428_/S vssd1 vssd1 vccd1 vccd1 _25380_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27110_ _27110_/CLK _27110_/D vssd1 vssd1 vccd1 vccd1 _27110_/Q sky130_fd_sc_hd__dfxtp_1
X_21534_ _21550_/A vssd1 vssd1 vccd1 vccd1 _21534_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24322_ _27545_/Q _24328_/B vssd1 vssd1 vccd1 vccd1 _24323_/A sky130_fd_sc_hd__and2_1
XFILLER_138_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24253_ _24253_/A _24287_/B vssd1 vssd1 vccd1 vccd1 _24254_/A sky130_fd_sc_hd__and2_1
X_27041_ _22948_/X _27041_/D vssd1 vssd1 vccd1 vccd1 _27041_/Q sky130_fd_sc_hd__dfxtp_1
X_21465_ _21459_/X _21460_/X _21461_/X _21462_/X _21463_/X _21464_/X vssd1 vssd1 vccd1
+ vccd1 _21466_/A sky130_fd_sc_hd__mux4_1
XFILLER_193_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23204_ _17453_/X _27139_/Q _23204_/S vssd1 vssd1 vccd1 vccd1 _23205_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20416_ _20408_/X _20409_/X _20410_/X _20411_/X _20412_/X _20413_/X vssd1 vssd1 vccd1
+ vccd1 _20417_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24184_ _27468_/Q _24184_/B vssd1 vssd1 vccd1 vccd1 _24185_/A sky130_fd_sc_hd__and2_1
XFILLER_179_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21396_ _21464_/A vssd1 vssd1 vccd1 vccd1 _21396_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23135_ _27108_/Q _17708_/X _23143_/S vssd1 vssd1 vccd1 vccd1 _23136_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20347_ _20347_/A vssd1 vssd1 vccd1 vccd1 _20347_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23066_ _27078_/Q _17715_/X _23070_/S vssd1 vssd1 vccd1 vccd1 _23067_/A sky130_fd_sc_hd__mux2_1
X_27943_ _27943_/A _15934_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20278_ _20267_/X _20269_/X _20271_/X _20273_/X _20274_/X _20275_/X vssd1 vssd1 vccd1
+ vccd1 _20279_/A sky130_fd_sc_hd__mux4_1
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22017_ _22017_/A vssd1 vssd1 vccd1 vccd1 _22084_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26825_ _22204_/X _26825_/D vssd1 vssd1 vccd1 vccd1 _26825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26756_ _21958_/X _26756_/D vssd1 vssd1 vccd1 vccd1 _26756_/Q sky130_fd_sc_hd__dfxtp_1
X_14770_ _14769_/X _26535_/Q _14773_/S vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23968_ _27848_/Q _27152_/Q _25897_/Q _25865_/Q _23967_/X _23944_/X vssd1 vssd1 vccd1
+ vccd1 _23968_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13721_ _13902_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13721_/Y sky130_fd_sc_hd__nor2_1
X_25707_ _25723_/A vssd1 vssd1 vccd1 vccd1 _25707_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22919_ _22907_/X _22908_/X _22909_/X _22910_/X _22911_/X _22912_/X vssd1 vssd1 vccd1
+ vccd1 _22920_/A sky130_fd_sc_hd__mux4_1
X_26687_ _21716_/X _26687_/D vssd1 vssd1 vccd1 vccd1 _26687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23899_ _23946_/A vssd1 vssd1 vccd1 vccd1 _23899_/X sky130_fd_sc_hd__buf_2
XFILLER_186_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16440_ _16779_/A _16440_/B vssd1 vssd1 vccd1 vccd1 _16441_/B sky130_fd_sc_hd__xor2_1
XFILLER_186_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13652_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25638_ _25638_/A vssd1 vssd1 vccd1 vccd1 _25638_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16744_/A _16371_/B vssd1 vssd1 vccd1 vccd1 _16396_/B sky130_fd_sc_hd__xor2_1
X_13583_ _13940_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13583_/Y sky130_fd_sc_hd__nor2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25569_ _25569_/A vssd1 vssd1 vccd1 vccd1 _25569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18110_ _18412_/A vssd1 vssd1 vccd1 vccd1 _18110_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15322_ _26303_/Q _13405_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15323_/A sky130_fd_sc_hd__mux2_1
X_27308_ _27308_/CLK _27308_/D vssd1 vssd1 vccd1 vccd1 _27308_/Q sky130_fd_sc_hd__dfxtp_1
X_19090_ _18996_/X _19088_/X _19089_/X vssd1 vssd1 vccd1 vccd1 _19090_/X sky130_fd_sc_hd__o21a_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18041_ _18182_/A vssd1 vssd1 vccd1 vccd1 _18041_/X sky130_fd_sc_hd__clkbuf_2
X_15253_ _15253_/A vssd1 vssd1 vccd1 vccd1 _26334_/D sky130_fd_sc_hd__clkbuf_1
X_27239_ _27263_/CLK _27239_/D vssd1 vssd1 vccd1 vccd1 _27239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14204_ _26727_/Q _14199_/X _14194_/X _14203_/Y vssd1 vssd1 vccd1 vccd1 _26727_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15184_ _26364_/Q _13414_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _26752_/Q _14130_/X _14133_/X _14134_/Y vssd1 vssd1 vccd1 vccd1 _26752_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19992_ _25639_/A vssd1 vssd1 vccd1 vccd1 _20338_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14066_ _14331_/A _14070_/B vssd1 vssd1 vccd1 vccd1 _14066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18943_ _26942_/Q _26910_/Q _26878_/Q _26846_/Q _18875_/X _18790_/X vssd1 vssd1 vccd1
+ vccd1 _18943_/X sky130_fd_sc_hd__mux4_2
X_13017_ _13017_/A vssd1 vssd1 vccd1 vccd1 _13061_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18874_ _18775_/X _18873_/X _18785_/X vssd1 vssd1 vccd1 vccd1 _18874_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17825_ _26138_/Q _26074_/Q _27002_/Q _26970_/Q _17821_/X _17824_/X vssd1 vssd1 vccd1
+ vccd1 _17828_/A sky130_fd_sc_hd__mux4_1
XFILLER_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17756_ _27433_/Q vssd1 vssd1 vccd1 vccd1 _17756_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14968_ _14975_/A vssd1 vssd1 vccd1 vccd1 _15023_/A sky130_fd_sc_hd__clkbuf_2
X_16707_ _16708_/A _16708_/B vssd1 vssd1 vccd1 vccd1 _16707_/Y sky130_fd_sc_hd__nor2_1
X_13919_ _13919_/A vssd1 vssd1 vccd1 vccd1 _13919_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17687_ _25915_/Q _17686_/X _17690_/S vssd1 vssd1 vccd1 vccd1 _17688_/A sky130_fd_sc_hd__mux2_1
X_14899_ _14727_/X _26484_/Q _14907_/S vssd1 vssd1 vccd1 vccd1 _14900_/A sky130_fd_sc_hd__mux2_1
X_19426_ _19471_/A _19426_/B _19426_/C vssd1 vssd1 vccd1 vccd1 _19427_/A sky130_fd_sc_hd__and3_1
X_16638_ _16638_/A _16638_/B vssd1 vssd1 vccd1 vccd1 _16638_/X sky130_fd_sc_hd__or2_1
XFILLER_63_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19357_ _26543_/Q _26511_/Q _26479_/Q _27055_/Q _19242_/X _19287_/X vssd1 vssd1 vccd1
+ vccd1 _19357_/X sky130_fd_sc_hd__mux4_1
X_16569_ _16569_/A vssd1 vssd1 vccd1 vccd1 _16888_/B sky130_fd_sc_hd__inv_2
XFILLER_200_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18308_ _18300_/X _18303_/X _18307_/X _18285_/X _18238_/X vssd1 vssd1 vccd1 vccd1
+ _18309_/C sky130_fd_sc_hd__a221o_1
X_19288_ _26540_/Q _26508_/Q _26476_/Q _27052_/Q _19242_/X _19287_/X vssd1 vssd1 vccd1
+ vccd1 _19288_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18239_ _18230_/X _18232_/X _18237_/X _18168_/X _18238_/X vssd1 vssd1 vccd1 vccd1
+ _18240_/C sky130_fd_sc_hd__a221o_1
XFILLER_198_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21250_ _21250_/A vssd1 vssd1 vccd1 vccd1 _21250_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20201_ _20249_/A vssd1 vssd1 vccd1 vccd1 _20201_/X sky130_fd_sc_hd__clkbuf_1
X_21181_ _21213_/A vssd1 vssd1 vccd1 vccd1 _21181_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20132_ _20164_/A vssd1 vssd1 vccd1 vccd1 _20132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20063_ _20079_/A vssd1 vssd1 vccd1 vccd1 _20063_/X sky130_fd_sc_hd__clkbuf_1
X_24940_ _24940_/A vssd1 vssd1 vccd1 vccd1 _24962_/A sky130_fd_sc_hd__clkbuf_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24871_ _27650_/Q _24861_/X _24870_/Y _24864_/X vssd1 vssd1 vccd1 vccd1 _27650_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater240 _27744_/CLK vssd1 vssd1 vccd1 vccd1 _27745_/CLK sky130_fd_sc_hd__clkbuf_1
X_26610_ _21450_/X _26610_/D vssd1 vssd1 vccd1 vccd1 _26610_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater251 _27536_/CLK vssd1 vssd1 vccd1 vccd1 _27604_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater262 _27172_/CLK vssd1 vssd1 vccd1 vccd1 _27536_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23822_ _23820_/X _23821_/X _23846_/S vssd1 vssd1 vccd1 vccd1 _23822_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27590_ _27592_/CLK _27590_/D vssd1 vssd1 vccd1 vccd1 _27590_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater273 _27475_/CLK vssd1 vssd1 vccd1 vccd1 _27600_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater284 _27484_/CLK vssd1 vssd1 vccd1 vccd1 _27520_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _18032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater295 _27245_/CLK vssd1 vssd1 vccd1 vccd1 _27262_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_318 _18973_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26541_ _21204_/X _26541_/D vssd1 vssd1 vccd1 vccd1 _26541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23753_ _23745_/X _23750_/X _23795_/S vssd1 vssd1 vccd1 vccd1 _23753_/X sky130_fd_sc_hd__mux2_1
X_20965_ _20953_/X _20954_/X _20955_/X _20956_/X _20958_/X _20960_/X vssd1 vssd1 vccd1
+ vccd1 _20966_/A sky130_fd_sc_hd__mux4_1
XANTENNA_329 _24005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22704_ _22772_/A vssd1 vssd1 vccd1 vccd1 _22704_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26472_ _20966_/X _26472_/D vssd1 vssd1 vccd1 vccd1 _26472_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _20896_/A vssd1 vssd1 vccd1 vccd1 _20896_/X sky130_fd_sc_hd__clkbuf_1
X_23684_ _23684_/A vssd1 vssd1 vccd1 vccd1 _27247_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25423_ _25423_/A vssd1 vssd1 vccd1 vccd1 _27749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22635_ _22893_/A vssd1 vssd1 vccd1 vccd1 _22700_/A sky130_fd_sc_hd__buf_2
XFILLER_55_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22566_ _22598_/A vssd1 vssd1 vccd1 vccd1 _22566_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25354_ _25354_/A _27518_/Q vssd1 vssd1 vccd1 vccd1 _25355_/B sky130_fd_sc_hd__xor2_1
XFILLER_107_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21517_ _21549_/A vssd1 vssd1 vccd1 vccd1 _21517_/X sky130_fd_sc_hd__clkbuf_2
X_24305_ _24305_/A _24384_/B vssd1 vssd1 vccd1 vccd1 _27434_/D sky130_fd_sc_hd__nor2_1
XFILLER_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22497_ _22487_/X _22488_/X _22489_/X _22490_/X _22491_/X _22492_/X vssd1 vssd1 vccd1
+ vccd1 _22498_/A sky130_fd_sc_hd__mux4_1
XFILLER_142_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25285_ _27539_/Q _27509_/Q vssd1 vssd1 vccd1 vccd1 _25287_/A sky130_fd_sc_hd__or2_1
XFILLER_103_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27024_ _22886_/X _27024_/D vssd1 vssd1 vccd1 vccd1 _27024_/Q sky130_fd_sc_hd__dfxtp_1
X_21448_ _21464_/A vssd1 vssd1 vccd1 vccd1 _21448_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24236_ _24304_/A vssd1 vssd1 vccd1 vccd1 _24256_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24167_ _27460_/Q _24173_/B vssd1 vssd1 vccd1 vccd1 _24168_/A sky130_fd_sc_hd__and2_1
X_21379_ _21373_/X _21374_/X _21375_/X _21376_/X _21377_/X _21378_/X vssd1 vssd1 vccd1
+ vccd1 _21380_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23118_ _23118_/A vssd1 vssd1 vccd1 vccd1 _27100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24098_ _27397_/Q _24106_/B vssd1 vssd1 vccd1 vccd1 _24099_/A sky130_fd_sc_hd__and2_1
XFILLER_27_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27926_ _27926_/A _15960_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
X_15940_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15940_/Y sky130_fd_sc_hd__inv_2
X_23049_ _23049_/A vssd1 vssd1 vccd1 vccd1 _27070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27857_ _27857_/CLK _27857_/D vssd1 vssd1 vccd1 vccd1 _27857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15871_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15871_/Y sky130_fd_sc_hd__inv_2
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17610_ _17434_/X _25878_/Q _17612_/S vssd1 vssd1 vccd1 vccd1 _17611_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26808_ _22138_/X _26808_/D vssd1 vssd1 vccd1 vccd1 _26808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14822_ _26518_/Q _13331_/X _14824_/S vssd1 vssd1 vccd1 vccd1 _14823_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _27688_/Q vssd1 vssd1 vccd1 vccd1 _25543_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27788_ _27788_/CLK _27788_/D vssd1 vssd1 vccd1 vccd1 _27788_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17541_ _17541_/A vssd1 vssd1 vccd1 vccd1 _25847_/D sky130_fd_sc_hd__clkbuf_1
X_26739_ _21894_/X _26739_/D vssd1 vssd1 vccd1 vccd1 _26739_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14753_/A vssd1 vssd1 vccd1 vccd1 _14753_/X sky130_fd_sc_hd__buf_2
XFILLER_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _26896_/Q _13697_/X _13692_/X _13703_/Y vssd1 vssd1 vccd1 vccd1 _26896_/D
+ sky130_fd_sc_hd__a31o_1
X_17472_ _27423_/Q vssd1 vssd1 vccd1 vccd1 _17472_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14684_ _25106_/A vssd1 vssd1 vccd1 vccd1 _14988_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19211_ _19209_/X _19210_/X _19211_/S vssd1 vssd1 vccd1 vccd1 _19211_/X sky130_fd_sc_hd__mux2_1
X_16423_ _16428_/A _16359_/A _16447_/C _16447_/D _16369_/A vssd1 vssd1 vccd1 vccd1
+ _16424_/B sky130_fd_sc_hd__o41a_1
X_13635_ _26920_/Q _13626_/X _13629_/X _13634_/Y vssd1 vssd1 vccd1 vccd1 _26920_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19142_ _26150_/Q _26086_/Q _27014_/Q _26982_/Q _19049_/X _19070_/X vssd1 vssd1 vccd1
+ vccd1 _19143_/B sky130_fd_sc_hd__mux4_1
X_16354_ _17674_/B _16508_/B vssd1 vssd1 vccd1 vccd1 _16354_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13566_ _26942_/Q _13558_/X _13553_/X _13565_/Y vssd1 vssd1 vccd1 vccd1 _26942_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ _15305_/A vssd1 vssd1 vccd1 vccd1 _26311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19073_ _19485_/A vssd1 vssd1 vccd1 vccd1 _19073_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16285_ _16109_/A _24297_/A _16593_/A vssd1 vssd1 vccd1 vccd1 _16801_/A sky130_fd_sc_hd__o21ai_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13497_ _16277_/A vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18024_ _26400_/Q _26368_/Q _26336_/Q _26304_/Q _17877_/X _17943_/X vssd1 vssd1 vccd1
+ vccd1 _18024_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15236_ _15247_/A vssd1 vssd1 vccd1 vccd1 _15245_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _26372_/Q _13389_/X _15173_/S vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14118_ _14383_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14118_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15098_ _15098_/A vssd1 vssd1 vccd1 vccd1 _26403_/D sky130_fd_sc_hd__clkbuf_1
X_19975_ _19991_/A vssd1 vssd1 vccd1 vccd1 _19975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14049_ _14521_/A vssd1 vssd1 vccd1 vccd1 _14406_/A sky130_fd_sc_hd__clkbuf_2
X_18926_ _18926_/A vssd1 vssd1 vccd1 vccd1 _24398_/A sky130_fd_sc_hd__buf_4
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18857_ _26139_/Q _26075_/Q _27003_/Q _26971_/Q _18807_/X _18810_/X vssd1 vssd1 vccd1
+ vccd1 _18858_/B sky130_fd_sc_hd__mux4_1
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17808_ _18177_/A vssd1 vssd1 vccd1 vccd1 _18387_/A sky130_fd_sc_hd__buf_4
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18788_ _19208_/A vssd1 vssd1 vccd1 vccd1 _18788_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _17739_/A vssd1 vssd1 vccd1 vccd1 _25931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20750_ _20738_/X _20739_/X _20740_/X _20741_/X _20742_/X _20743_/X vssd1 vssd1 vccd1
+ vccd1 _20751_/A sky130_fd_sc_hd__mux4_1
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19409_ _19409_/A _19409_/B vssd1 vssd1 vccd1 vccd1 _19409_/X sky130_fd_sc_hd__or2_1
X_20681_ _20681_/A vssd1 vssd1 vccd1 vccd1 _20681_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22420_ _22436_/A vssd1 vssd1 vccd1 vccd1 _22420_/X sky130_fd_sc_hd__clkbuf_1
X_22351_ _22523_/A vssd1 vssd1 vccd1 vccd1 _22421_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21302_ _21302_/A vssd1 vssd1 vccd1 vccd1 _21302_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25070_ _27230_/Q vssd1 vssd1 vccd1 vccd1 _25070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22282_ _22348_/A vssd1 vssd1 vccd1 vccd1 _22282_/X sky130_fd_sc_hd__clkbuf_1
X_24021_ _23990_/X _24019_/X _24020_/X _24005_/X vssd1 vssd1 vccd1 vccd1 _27298_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21233_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21164_ _21212_/A vssd1 vssd1 vccd1 vccd1 _21164_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20115_ _20163_/A vssd1 vssd1 vccd1 vccd1 _20115_/X sky130_fd_sc_hd__clkbuf_1
X_25972_ _26069_/CLK _25972_/D vssd1 vssd1 vccd1 vccd1 _25972_/Q sky130_fd_sc_hd__dfxtp_1
X_21095_ _21127_/A vssd1 vssd1 vccd1 vccd1 _21095_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27711_ _27711_/CLK _27711_/D vssd1 vssd1 vccd1 vccd1 _27711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20046_ _20078_/A vssd1 vssd1 vccd1 vccd1 _20046_/X sky130_fd_sc_hd__clkbuf_1
X_24923_ _24937_/A _24923_/B vssd1 vssd1 vccd1 vccd1 _24923_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27642_ _27642_/CLK _27642_/D vssd1 vssd1 vccd1 vccd1 _27642_/Q sky130_fd_sc_hd__dfxtp_1
X_24854_ _24863_/A _24854_/B vssd1 vssd1 vccd1 vccd1 _24854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23805_ _25917_/Q _25983_/Q _25816_/Q _26015_/Q _23804_/X _23786_/X vssd1 vssd1 vccd1
+ vccd1 _23805_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27573_ _27573_/CLK _27573_/D vssd1 vssd1 vccd1 vccd1 _27573_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_104 _19447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _22540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24785_ _24861_/A vssd1 vssd1 vccd1 vccd1 _24785_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _21997_/A vssd1 vssd1 vccd1 vccd1 _21997_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_126 _22616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 _23598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26524_ _21142_/X _26524_/D vssd1 vssd1 vccd1 vccd1 _26524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _13116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23736_ _27374_/Q _24050_/B vssd1 vssd1 vccd1 vccd1 _23737_/A sky130_fd_sc_hd__and2_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20948_/A vssd1 vssd1 vccd1 vccd1 _20948_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_159 _13382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26455_ _20912_/X _26455_/D vssd1 vssd1 vccd1 vccd1 _26455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23667_ _23667_/A vssd1 vssd1 vccd1 vccd1 _27239_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20879_ _20864_/X _20865_/X _20866_/X _20867_/X _20870_/X _20874_/X vssd1 vssd1 vccd1
+ vccd1 _20880_/A sky130_fd_sc_hd__mux4_1
XFILLER_201_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25406_ _25406_/A vssd1 vssd1 vccd1 vccd1 _27741_/D sky130_fd_sc_hd__clkbuf_1
X_13420_ _14810_/A vssd1 vssd1 vccd1 vccd1 _13420_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_197_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22618_ _22686_/A vssd1 vssd1 vccd1 vccd1 _22618_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26386_ _20661_/X _26386_/D vssd1 vssd1 vccd1 vccd1 _26386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23598_ _23598_/A vssd1 vssd1 vccd1 vccd1 _23617_/A sky130_fd_sc_hd__clkbuf_1
X_25337_ _27717_/Q _25308_/X _25336_/Y _13423_/X vssd1 vssd1 vccd1 vccd1 _27717_/D
+ sky130_fd_sc_hd__o211a_1
X_13351_ _26992_/Q _13350_/X _13351_/S vssd1 vssd1 vccd1 vccd1 _13352_/A sky130_fd_sc_hd__mux2_1
X_22549_ _22597_/A vssd1 vssd1 vccd1 vccd1 _22549_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16070_ _16402_/A vssd1 vssd1 vccd1 vccd1 _16094_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25268_ _25241_/B _25250_/X _25265_/Y _25267_/Y _25258_/B vssd1 vssd1 vccd1 vccd1
+ _25272_/B sky130_fd_sc_hd__a311oi_4
X_13282_ _13304_/A vssd1 vssd1 vccd1 vccd1 _13291_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15021_ _15758_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _15021_/Y sky130_fd_sc_hd__nor2_1
X_27007_ _22832_/X _27007_/D vssd1 vssd1 vccd1 vccd1 _27007_/Q sky130_fd_sc_hd__dfxtp_1
X_24219_ _25615_/A _24222_/B vssd1 vssd1 vccd1 vccd1 _27378_/D sky130_fd_sc_hd__nor2_1
XFILLER_163_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25199_ _25221_/A _25199_/B vssd1 vssd1 vccd1 vccd1 _25199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19760_ _19745_/X _19747_/X _19749_/X _19751_/X _19752_/X _19753_/X vssd1 vssd1 vccd1
+ vccd1 _19761_/A sky130_fd_sc_hd__mux4_1
X_16972_ _16979_/A _24636_/A _16982_/C _16982_/D vssd1 vssd1 vccd1 vccd1 _16973_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_150_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15923_ _15924_/A vssd1 vssd1 vccd1 vccd1 _15923_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18711_ _26018_/Q _17702_/X _18713_/S vssd1 vssd1 vccd1 vccd1 _18712_/A sky130_fd_sc_hd__mux2_1
X_19691_ _19691_/A vssd1 vssd1 vccd1 vccd1 _19691_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18642_ _18642_/A vssd1 vssd1 vccd1 vccd1 _25987_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15854_ _15854_/A vssd1 vssd1 vccd1 vccd1 _26074_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_842 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14805_ _14804_/X _26524_/Q _14805_/S vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__mux2_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _18468_/X _18568_/X _18572_/X _18016_/X vssd1 vssd1 vccd1 vccd1 _18582_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15785_ _15853_/S vssd1 vssd1 vccd1 vccd1 _15794_/S sky130_fd_sc_hd__clkbuf_2
X_12997_ _12997_/A vssd1 vssd1 vccd1 vccd1 _27800_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _17523_/X _25842_/Q _17524_/S vssd1 vssd1 vccd1 vccd1 _17525_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _14736_/A vssd1 vssd1 vccd1 vccd1 _26546_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _17455_/A vssd1 vssd1 vccd1 vccd1 _25820_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _15741_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14667_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16406_ _16406_/A vssd1 vssd1 vccd1 vccd1 _16774_/A sky130_fd_sc_hd__clkbuf_2
X_13618_ _26927_/Q _13613_/X _13616_/X _13617_/Y vssd1 vssd1 vccd1 vccd1 _26927_/D
+ sky130_fd_sc_hd__a31o_1
X_17386_ _17384_/X _17385_/X _17386_/S vssd1 vssd1 vccd1 vccd1 _17386_/X sky130_fd_sc_hd__mux2_2
X_14598_ _26595_/Q _14589_/X _14592_/X _14597_/Y vssd1 vssd1 vccd1 vccd1 _26595_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19125_ _19073_/X _19124_/X _19076_/X vssd1 vssd1 vccd1 vccd1 _19125_/X sky130_fd_sc_hd__o21a_1
X_16337_ _16753_/B _16349_/B vssd1 vssd1 vccd1 vccd1 _16337_/X sky130_fd_sc_hd__or2_1
XFILLER_173_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _27342_/Q _13063_/X _13064_/X _27310_/Q _13196_/X vssd1 vssd1 vccd1 vccd1
+ _14507_/A sky130_fd_sc_hd__a221oi_4
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19056_ _26530_/Q _26498_/Q _26466_/Q _27042_/Q _18984_/X _19032_/X vssd1 vssd1 vccd1
+ vccd1 _19056_/X sky130_fd_sc_hd__mux4_1
X_16268_ _26059_/Q _16274_/B _16274_/C vssd1 vssd1 vccd1 vccd1 _16268_/X sky130_fd_sc_hd__and3_1
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18007_ _18479_/A vssd1 vssd1 vccd1 vccd1 _24392_/A sky130_fd_sc_hd__clkbuf_4
X_15219_ _14750_/X _26349_/Q _15223_/S vssd1 vssd1 vccd1 vccd1 _15220_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16199_ _16172_/X _16194_/X _16196_/Y _16197_/X _16198_/X vssd1 vssd1 vccd1 vccd1
+ _16326_/A sky130_fd_sc_hd__o41a_1
XFILLER_160_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19958_ _19990_/A vssd1 vssd1 vccd1 vccd1 _19958_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18909_ _19486_/A vssd1 vssd1 vccd1 vccd1 _18909_/X sky130_fd_sc_hd__buf_2
X_19889_ _19889_/A vssd1 vssd1 vccd1 vccd1 _19889_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21920_ _21920_/A vssd1 vssd1 vccd1 vccd1 _21920_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21851_ _21899_/A vssd1 vssd1 vccd1 vccd1 _21851_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20802_ _21149_/A vssd1 vssd1 vccd1 vccd1 _20867_/A sky130_fd_sc_hd__clkbuf_2
X_21782_ _21814_/A vssd1 vssd1 vccd1 vccd1 _21782_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24570_ _27646_/Q _24576_/B vssd1 vssd1 vccd1 vccd1 _24571_/A sky130_fd_sc_hd__and2_1
XFILLER_64_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23521_ _24835_/B _27198_/Q _23525_/S vssd1 vssd1 vccd1 vccd1 _23522_/B sky130_fd_sc_hd__mux2_1
XFILLER_196_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20733_ _20733_/A vssd1 vssd1 vccd1 vccd1 _20733_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26240_ _20153_/X _26240_/D vssd1 vssd1 vccd1 vccd1 _26240_/Q sky130_fd_sc_hd__dfxtp_1
X_23452_ input12/X _23442_/X _23451_/X _23447_/X vssd1 vssd1 vccd1 vccd1 _27174_/D
+ sky130_fd_sc_hd__o211a_1
X_20664_ _20652_/X _20653_/X _20654_/X _20655_/X _20656_/X _20657_/X vssd1 vssd1 vccd1
+ vccd1 _20665_/A sky130_fd_sc_hd__mux4_1
XFILLER_91_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22403_ _22435_/A vssd1 vssd1 vccd1 vccd1 _22403_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23383_ _27242_/Q vssd1 vssd1 vccd1 vccd1 _23383_/Y sky130_fd_sc_hd__inv_2
X_26171_ _19909_/X _26171_/D vssd1 vssd1 vccd1 vccd1 _26171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20595_ _20595_/A vssd1 vssd1 vccd1 vccd1 _20595_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25122_ _25122_/A _25122_/B vssd1 vssd1 vccd1 vccd1 _25123_/B sky130_fd_sc_hd__xnor2_1
X_22334_ _22350_/A vssd1 vssd1 vccd1 vccd1 _22334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22265_ _22523_/A vssd1 vssd1 vccd1 vccd1 _22335_/A sky130_fd_sc_hd__clkbuf_2
X_25053_ _25921_/Q _25987_/Q _25820_/Q _26019_/Q _25052_/X _25027_/X vssd1 vssd1 vccd1
+ vccd1 _25053_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24004_ _27091_/Q _24001_/X _24002_/X _27123_/Q _24003_/X vssd1 vssd1 vccd1 vccd1
+ _24004_/X sky130_fd_sc_hd__a221o_1
XFILLER_133_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21216_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21216_/X sky130_fd_sc_hd__clkbuf_2
X_22196_ _22262_/A vssd1 vssd1 vccd1 vccd1 _22196_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21147_ _21147_/A vssd1 vssd1 vccd1 vccd1 _21213_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21078_ _21126_/A vssd1 vssd1 vccd1 vccd1 _21078_/X sky130_fd_sc_hd__clkbuf_1
X_25955_ _27327_/CLK _25955_/D vssd1 vssd1 vccd1 vccd1 _25955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12920_ input57/X input58/X input59/X input60/X vssd1 vssd1 vccd1 vccd1 _12921_/B
+ sky130_fd_sc_hd__and4_1
X_24906_ _24906_/A _24910_/C vssd1 vssd1 vccd1 vccd1 _24907_/B sky130_fd_sc_hd__xnor2_1
X_20029_ _20077_/A vssd1 vssd1 vccd1 vccd1 _20029_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25886_ _27141_/CLK _25886_/D vssd1 vssd1 vccd1 vccd1 _25886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27625_ _27625_/CLK _27625_/D vssd1 vssd1 vccd1 vccd1 _27625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24837_ _24844_/B _24837_/B vssd1 vssd1 vccd1 vccd1 _24838_/B sky130_fd_sc_hd__or2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27556_ _27558_/CLK _27556_/D vssd1 vssd1 vccd1 vccd1 _27556_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15570_/A vssd1 vssd1 vccd1 vccd1 _26194_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24768_ _27621_/Q _24758_/X _24767_/Y _24760_/X vssd1 vssd1 vccd1 vccd1 _27621_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14521_ _14521_/A vssd1 vssd1 vccd1 vccd1 _15775_/A sky130_fd_sc_hd__clkbuf_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26507_ _21088_/X _26507_/D vssd1 vssd1 vccd1 vccd1 _26507_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23719_ _23719_/A vssd1 vssd1 vccd1 vccd1 _27263_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27487_ _27488_/CLK _27487_/D vssd1 vssd1 vccd1 vccd1 _27487_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24699_ _24396_/A _24687_/X _24698_/X _24690_/X vssd1 vssd1 vccd1 vccd1 _27597_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _25931_/Q _25997_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17241_/B sky130_fd_sc_hd__mux2_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14452_/A vssd1 vssd1 vccd1 vccd1 _15725_/A sky130_fd_sc_hd__clkbuf_2
X_26438_ _20845_/X _26438_/D vssd1 vssd1 vccd1 vccd1 _26438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ _26976_/Q _13401_/X _13415_/S vssd1 vssd1 vccd1 vccd1 _13404_/A sky130_fd_sc_hd__mux2_1
X_17171_ _17120_/X _17170_/X _17159_/X vssd1 vssd1 vccd1 vccd1 _17171_/X sky130_fd_sc_hd__a21bo_1
X_14383_ _14383_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _14383_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26369_ _20597_/X _26369_/D vssd1 vssd1 vccd1 vccd1 _26369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16122_ _27406_/Q _16144_/B vssd1 vssd1 vccd1 vccd1 _16122_/Y sky130_fd_sc_hd__nand2_1
X_13334_ _14724_/A vssd1 vssd1 vccd1 vccd1 _13334_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ _27476_/Q vssd1 vssd1 vccd1 vccd1 _16053_/Y sky130_fd_sc_hd__inv_2
X_13265_ _27026_/Q _13099_/X _13269_/S vssd1 vssd1 vccd1 vccd1 _13266_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15004_ _15741_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ _27278_/Q _13237_/B vssd1 vssd1 vccd1 vccd1 _13196_/X sky130_fd_sc_hd__and2_2
XFILLER_97_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19812_ _19812_/A vssd1 vssd1 vccd1 vccd1 _19812_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19743_ _19743_/A vssd1 vssd1 vccd1 vccd1 _19743_/X sky130_fd_sc_hd__clkbuf_1
X_16955_ _27581_/Q _27580_/Q _27579_/Q _27578_/Q vssd1 vssd1 vccd1 vccd1 _24626_/D
+ sky130_fd_sc_hd__or4bb_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15906_ _15906_/A vssd1 vssd1 vccd1 vccd1 _15906_/Y sky130_fd_sc_hd__inv_2
X_16886_ _16884_/X _16801_/X _16885_/X _16877_/X vssd1 vssd1 vccd1 vccd1 _24249_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_19674_ _19659_/X _19661_/X _19663_/X _19665_/X _19666_/X _19667_/X vssd1 vssd1 vccd1
+ vccd1 _19675_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18625_ _18625_/A vssd1 vssd1 vccd1 vccd1 _25979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15837_ _15837_/A vssd1 vssd1 vccd1 vccd1 _26082_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15768_ _26112_/Q _15760_/X _15766_/X _15767_/Y vssd1 vssd1 vccd1 vccd1 _26112_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18556_ _26168_/Q _26104_/Q _27032_/Q _27000_/Q _18455_/X _18011_/X vssd1 vssd1 vccd1
+ vccd1 _18557_/A sky130_fd_sc_hd__mux4_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17507_ _17507_/A vssd1 vssd1 vccd1 vccd1 _25836_/D sky130_fd_sc_hd__clkbuf_1
X_14719_ _14718_/X _26551_/Q _14725_/S vssd1 vssd1 vccd1 vccd1 _14720_/A sky130_fd_sc_hd__mux2_1
X_18487_ _26420_/Q _26388_/Q _26356_/Q _26324_/Q _18462_/X _18486_/X vssd1 vssd1 vccd1
+ vccd1 _18487_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15699_ _15699_/A _15703_/B vssd1 vssd1 vccd1 vccd1 _15699_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17438_ _17437_/X _25815_/Q _17438_/S vssd1 vssd1 vccd1 vccd1 _17439_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_15 _25989_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_26 _27142_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_37 _18481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 _18001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17369_ _27856_/Q _27160_/Q _25905_/Q _25873_/Q _17325_/X _17181_/A vssd1 vssd1 vccd1
+ vccd1 _17369_/X sky130_fd_sc_hd__mux4_1
XFILLER_146_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_59 _18251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19108_ _19108_/A vssd1 vssd1 vccd1 vccd1 _26052_/D sky130_fd_sc_hd__clkbuf_1
X_20380_ _20412_/A vssd1 vssd1 vccd1 vccd1 _20380_/X sky130_fd_sc_hd__clkbuf_2
X_19039_ _19338_/A vssd1 vssd1 vccd1 vccd1 _19039_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22050_ _22050_/A vssd1 vssd1 vccd1 vccd1 _22050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21001_ _20991_/X _20992_/X _20993_/X _20994_/X _20995_/X _20996_/X vssd1 vssd1 vccd1
+ vccd1 _21002_/A sky130_fd_sc_hd__mux4_1
XFILLER_82_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25740_ _17428_/X _27827_/Q _25746_/S vssd1 vssd1 vccd1 vccd1 _25741_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22952_ _22952_/A vssd1 vssd1 vccd1 vccd1 _22952_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21903_ _21895_/X _21896_/X _21897_/X _21898_/X _21899_/X _21900_/X vssd1 vssd1 vccd1
+ vccd1 _21904_/A sky130_fd_sc_hd__mux4_1
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25671_ _25654_/X _25656_/X _25658_/X _25660_/X _25661_/X _25662_/X vssd1 vssd1 vccd1
+ vccd1 _25672_/A sky130_fd_sc_hd__mux4_1
X_22883_ _22869_/X _22870_/X _22871_/X _22872_/X _22874_/X _22876_/X vssd1 vssd1 vccd1
+ vccd1 _22884_/A sky130_fd_sc_hd__mux4_1
XFILLER_83_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27410_ _27410_/CLK _27410_/D vssd1 vssd1 vccd1 vccd1 _27410_/Q sky130_fd_sc_hd__dfxtp_1
X_24622_ _27670_/Q _24624_/B vssd1 vssd1 vccd1 vccd1 _24623_/A sky130_fd_sc_hd__and2_1
X_21834_ _21834_/A vssd1 vssd1 vccd1 vccd1 _21834_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27341_ _27341_/CLK _27341_/D vssd1 vssd1 vccd1 vccd1 _27341_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24553_ _24553_/A vssd1 vssd1 vccd1 vccd1 _27538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21765_ _21813_/A vssd1 vssd1 vccd1 vccd1 _21765_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_905 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23504_ _25625_/S vssd1 vssd1 vccd1 vccd1 _25430_/B sky130_fd_sc_hd__buf_2
XFILLER_93_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20716_ _20703_/X _20705_/X _20707_/X _20709_/X _20710_/X _20711_/X vssd1 vssd1 vccd1
+ vccd1 _20717_/A sky130_fd_sc_hd__mux4_1
X_27272_ _27411_/CLK _27272_/D vssd1 vssd1 vccd1 vccd1 _27272_/Q sky130_fd_sc_hd__dfxtp_1
X_24484_ _24484_/A vssd1 vssd1 vccd1 vccd1 _27517_/D sky130_fd_sc_hd__clkbuf_1
X_21696_ _21696_/A vssd1 vssd1 vccd1 vccd1 _21696_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_949 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26223_ _20091_/X _26223_/D vssd1 vssd1 vccd1 vccd1 _26223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23435_ _16998_/X _23429_/X _23433_/X _23434_/X vssd1 vssd1 vccd1 vccd1 _27167_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_196_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20647_ _20647_/A vssd1 vssd1 vccd1 vccd1 _20647_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26154_ _19849_/X _26154_/D vssd1 vssd1 vccd1 vccd1 _26154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20578_ _20566_/X _20567_/X _20568_/X _20569_/X _20570_/X _20571_/X vssd1 vssd1 vccd1
+ vccd1 _20579_/A sky130_fd_sc_hd__mux4_2
X_23366_ _27775_/Q vssd1 vssd1 vccd1 vccd1 _24792_/A sky130_fd_sc_hd__inv_2
XFILLER_178_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25105_ _25105_/A vssd1 vssd1 vccd1 vccd1 _27687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22317_ _22349_/A vssd1 vssd1 vccd1 vccd1 _22317_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26085_ _19612_/X _26085_/D vssd1 vssd1 vccd1 vccd1 _26085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23297_ _27740_/Q _23263_/Y _27735_/Q _23296_/Y vssd1 vssd1 vccd1 vccd1 _23297_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13050_ _13205_/A vssd1 vssd1 vccd1 vccd1 _13241_/S sky130_fd_sc_hd__clkbuf_4
X_25036_ _27833_/Q _27137_/Q _25882_/Q _25850_/Q _25018_/X _25035_/X vssd1 vssd1 vccd1
+ vccd1 _25036_/X sky130_fd_sc_hd__mux4_1
X_22248_ _22264_/A vssd1 vssd1 vccd1 vccd1 _22248_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22179_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26987_ _22762_/X _26987_/D vssd1 vssd1 vccd1 vccd1 _26987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16740_ _16747_/A _16742_/A _16739_/X vssd1 vssd1 vccd1 vccd1 _16740_/Y sky130_fd_sc_hd__o21ai_1
X_25938_ _27854_/CLK _25938_/D vssd1 vssd1 vccd1 vccd1 _25938_/Q sky130_fd_sc_hd__dfxtp_1
X_13952_ _26808_/Q _13949_/X _13944_/X _13951_/Y vssd1 vssd1 vccd1 vccd1 _26808_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16671_ _16700_/A _16700_/B _16500_/A vssd1 vssd1 vccd1 vccd1 _16672_/B sky130_fd_sc_hd__a21oi_1
XFILLER_19_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25869_ _27852_/CLK _25869_/D vssd1 vssd1 vccd1 vccd1 _25869_/Q sky130_fd_sc_hd__dfxtp_1
X_13883_ _26833_/Q _13880_/X _13873_/X _13882_/Y vssd1 vssd1 vccd1 vccd1 _26833_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18410_ _18410_/A _18317_/X vssd1 vssd1 vccd1 vccd1 _18410_/X sky130_fd_sc_hd__or2b_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15622_ _15622_/A vssd1 vssd1 vccd1 vccd1 _26170_/D sky130_fd_sc_hd__clkbuf_1
X_19390_ _27816_/Q _26577_/Q _26449_/Q _26129_/Q _19255_/X _19321_/X vssd1 vssd1 vccd1
+ vccd1 _19390_/X sky130_fd_sc_hd__mux4_1
X_27608_ _27608_/CLK _27608_/D vssd1 vssd1 vccd1 vccd1 _27608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18339_/X _18340_/X _18395_/A vssd1 vssd1 vccd1 vccd1 _18341_/X sky130_fd_sc_hd__mux2_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27539_ _27539_/CLK _27539_/D vssd1 vssd1 vccd1 vccd1 _27539_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15621_/S vssd1 vssd1 vccd1 vccd1 _15562_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14519_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _26827_/Q _26795_/Q _26763_/Q _26731_/Q _18175_/X _18199_/X vssd1 vssd1 vccd1
+ vccd1 _18272_/X sky130_fd_sc_hd__mux4_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _13058_/X _26232_/Q _15490_/S vssd1 vssd1 vccd1 vccd1 _15485_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17223_ _27083_/Q _27115_/Q _17234_/S vssd1 vssd1 vccd1 vccd1 _17223_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14435_ _26645_/Q _14421_/X _14416_/X _14434_/Y vssd1 vssd1 vccd1 vccd1 _26645_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 la1_data_in[13] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17154_ _27838_/Q _27142_/Q _25887_/Q _25855_/Q _17142_/X _17130_/X vssd1 vssd1 vccd1
+ vccd1 _17154_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput24 la1_data_in[23] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
X_14366_ _14393_/A vssd1 vssd1 vccd1 vccd1 _14376_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 la1_data_in[4] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput46 la1_oenb[14] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 la1_oenb[24] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
Xinput68 la1_oenb[5] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_4
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ _16486_/A vssd1 vssd1 vccd1 vccd1 _16106_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13317_ _27002_/Q _13240_/X _13317_/S vssd1 vssd1 vccd1 vccd1 _13318_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17085_ _17029_/X _17085_/B vssd1 vssd1 vccd1 vccd1 _17085_/X sky130_fd_sc_hd__and2b_1
X_14297_ _14311_/A vssd1 vssd1 vccd1 vccd1 _14297_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ _16266_/A vssd1 vssd1 vccd1 vccd1 _16036_/X sky130_fd_sc_hd__buf_2
X_13248_ _13304_/A vssd1 vssd1 vccd1 vccd1 _13317_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_184_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ _14779_/A vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__buf_2
XFILLER_42_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17987_ _26527_/Q _26495_/Q _26463_/Q _27039_/Q _17964_/X _17986_/X vssd1 vssd1 vccd1
+ vccd1 _17987_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19726_ _19726_/A vssd1 vssd1 vccd1 vccd1 _19726_/X sky130_fd_sc_hd__clkbuf_1
X_16938_ _18828_/A _24206_/A _24207_/A _27599_/Q vssd1 vssd1 vccd1 vccd1 _16945_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19657_ _19657_/A vssd1 vssd1 vccd1 vccd1 _19657_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _16755_/A _16753_/B _16868_/X vssd1 vssd1 vccd1 vccd1 _16869_/Y sky130_fd_sc_hd__o21ai_1
X_18608_ _24828_/A _18606_/X _24823_/A vssd1 vssd1 vccd1 vccd1 _18608_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19588_ _19588_/A vssd1 vssd1 vccd1 vccd1 _19588_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18539_ _18539_/A _18479_/X vssd1 vssd1 vccd1 vccd1 _18539_/X sky130_fd_sc_hd__or2b_1
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21550_ _21550_/A vssd1 vssd1 vccd1 vccd1 _21550_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20501_ _20501_/A vssd1 vssd1 vccd1 vccd1 _20501_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21481_ _21653_/A vssd1 vssd1 vccd1 vccd1 _21550_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23220_ _17476_/X _27146_/Q _23226_/S vssd1 vssd1 vccd1 vccd1 _23221_/A sky130_fd_sc_hd__mux2_1
X_20432_ _20776_/A vssd1 vssd1 vccd1 vccd1 _20501_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_146_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23151_ _23151_/A vssd1 vssd1 vccd1 vccd1 _27115_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20363_ _20427_/A vssd1 vssd1 vccd1 vccd1 _20363_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22102_ _22451_/A vssd1 vssd1 vccd1 vccd1 _22173_/A sky130_fd_sc_hd__clkbuf_2
X_23082_ _23082_/A vssd1 vssd1 vccd1 vccd1 _27085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20294_ _20286_/X _20287_/X _20288_/X _20289_/X _20290_/X _20291_/X vssd1 vssd1 vccd1
+ vccd1 _20295_/A sky130_fd_sc_hd__mux4_1
XFILLER_164_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22033_ _22016_/X _22018_/X _22020_/X _22022_/X _22023_/X _22024_/X vssd1 vssd1 vccd1
+ vccd1 _22034_/A sky130_fd_sc_hd__mux4_1
X_26910_ _22494_/X _26910_/D vssd1 vssd1 vccd1 vccd1 _26910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26841_ _22254_/X _26841_/D vssd1 vssd1 vccd1 vccd1 _26841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26772_ _22010_/X _26772_/D vssd1 vssd1 vccd1 vccd1 _26772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23984_ _25936_/Q _26002_/Q _25835_/Q _26034_/Q _23946_/X _23976_/X vssd1 vssd1 vccd1
+ vccd1 _23984_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25723_ _25723_/A vssd1 vssd1 vccd1 vccd1 _25723_/X sky130_fd_sc_hd__clkbuf_1
X_22935_ _22923_/X _22924_/X _22925_/X _22926_/X _22927_/X _22928_/X vssd1 vssd1 vccd1
+ vccd1 _22936_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25654_ _25721_/A vssd1 vssd1 vccd1 vccd1 _25654_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22866_ _22866_/A vssd1 vssd1 vccd1 vccd1 _22866_/X sky130_fd_sc_hd__clkbuf_1
X_24605_ _27662_/Q _24609_/B vssd1 vssd1 vccd1 vccd1 _24606_/A sky130_fd_sc_hd__and2_1
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21817_ _21809_/X _21810_/X _21811_/X _21812_/X _21813_/X _21814_/X vssd1 vssd1 vccd1
+ vccd1 _21818_/A sky130_fd_sc_hd__mux4_1
X_25585_ _25572_/X _25582_/X _25583_/X _24944_/B _25584_/X vssd1 vssd1 vccd1 vccd1
+ _25585_/X sky130_fd_sc_hd__o311a_1
XFILLER_145_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22797_ _22783_/X _22784_/X _22785_/X _22786_/X _22788_/X _22790_/X vssd1 vssd1 vccd1
+ vccd1 _22798_/A sky130_fd_sc_hd__mux4_1
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27324_ _27325_/CLK _27324_/D vssd1 vssd1 vccd1 vccd1 _27324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24536_ _24631_/A _24536_/B vssd1 vssd1 vccd1 vccd1 _24537_/A sky130_fd_sc_hd__and2_1
X_21748_ _21748_/A vssd1 vssd1 vccd1 vccd1 _21748_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_605 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27255_ _27778_/CLK _27255_/D vssd1 vssd1 vccd1 vccd1 _27255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24467_ _27631_/Q _24467_/B vssd1 vssd1 vccd1 vccd1 _24468_/A sky130_fd_sc_hd__and2_1
XFILLER_200_757 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21679_ _21667_/X _21670_/X _21673_/X _21676_/X _21677_/X _21678_/X vssd1 vssd1 vccd1
+ vccd1 _21680_/A sky130_fd_sc_hd__mux4_1
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _14220_/A vssd1 vssd1 vccd1 vccd1 _14220_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26206_ _20037_/X _26206_/D vssd1 vssd1 vccd1 vccd1 _26206_/Q sky130_fd_sc_hd__dfxtp_1
X_23418_ _23500_/B vssd1 vssd1 vccd1 vccd1 _23430_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_138_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27186_ _27589_/CLK _27186_/D vssd1 vssd1 vccd1 vccd1 _27186_/Q sky130_fd_sc_hd__dfxtp_1
X_24398_ _24398_/A _24400_/B vssd1 vssd1 vccd1 vccd1 _24399_/A sky130_fd_sc_hd__and2_1
XFILLER_153_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _14234_/B vssd1 vssd1 vccd1 vccd1 _14151_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26137_ _19791_/X _26137_/D vssd1 vssd1 vccd1 vccd1 _26137_/Q sky130_fd_sc_hd__dfxtp_1
X_23349_ _27773_/Q vssd1 vssd1 vccd1 vccd1 _24786_/A sky130_fd_sc_hd__inv_2
XFILLER_180_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _13102_/A vssd1 vssd1 vccd1 vccd1 _13102_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_153_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14082_ _26772_/Q _14076_/X _14080_/X _14081_/Y vssd1 vssd1 vccd1 vccd1 _26772_/D
+ sky130_fd_sc_hd__a31o_1
X_26068_ _26068_/CLK _26068_/D vssd1 vssd1 vccd1 vccd1 _26068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25019_ _27831_/Q _27135_/Q _25880_/Q _25848_/Q _25018_/X _24991_/X vssd1 vssd1 vccd1
+ vccd1 _25019_/X sky130_fd_sc_hd__mux4_1
X_13033_ _13201_/B vssd1 vssd1 vccd1 vccd1 _13176_/B sky130_fd_sc_hd__clkbuf_1
X_17910_ _18522_/S vssd1 vssd1 vccd1 vccd1 _17910_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18890_ _18888_/X _18889_/X _19539_/S vssd1 vssd1 vccd1 vccd1 _18890_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17841_ _18392_/A vssd1 vssd1 vccd1 vccd1 _17841_/X sky130_fd_sc_hd__buf_4
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17772_ _27438_/Q vssd1 vssd1 vccd1 vccd1 _17772_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14984_ _15723_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19511_ _19509_/X _19510_/X _19565_/S vssd1 vssd1 vccd1 vccd1 _19511_/X sky130_fd_sc_hd__mux2_1
X_13935_ _26813_/Q _13933_/X _13925_/X _13934_/Y vssd1 vssd1 vccd1 vccd1 _26813_/D
+ sky130_fd_sc_hd__a31o_1
X_16723_ _16084_/A _16721_/Y _16722_/X _16626_/A vssd1 vssd1 vccd1 vccd1 _16723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16654_ _16654_/A _16654_/B vssd1 vssd1 vccd1 vccd1 _16654_/Y sky130_fd_sc_hd__xnor2_1
X_19442_ _26291_/Q _26259_/Q _26227_/Q _26195_/Q _19441_/X _19352_/X vssd1 vssd1 vccd1
+ vccd1 _19442_/X sky130_fd_sc_hd__mux4_1
X_13866_ _13872_/A vssd1 vssd1 vccd1 vccd1 _13920_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15605_ _15605_/A vssd1 vssd1 vccd1 vccd1 _26178_/D sky130_fd_sc_hd__clkbuf_1
X_16585_ _16916_/A _16585_/B vssd1 vssd1 vccd1 vccd1 _16913_/B sky130_fd_sc_hd__nand2_1
X_19373_ _26416_/Q _26384_/Q _26352_/Q _26320_/Q _18900_/X _18901_/X vssd1 vssd1 vccd1
+ vccd1 _19373_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13797_ _13889_/A _13799_/B vssd1 vssd1 vccd1 vccd1 _13797_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18324_ _18324_/A vssd1 vssd1 vccd1 vccd1 _18324_/X sky130_fd_sc_hd__clkbuf_2
X_15536_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15545_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_188_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18255_ _26154_/Q _26090_/Q _27018_/Q _26986_/Q _18182_/X _18228_/X vssd1 vssd1 vccd1
+ vccd1 _18256_/A sky130_fd_sc_hd__mux4_1
XFILLER_72_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15467_ _26239_/Q _13405_/X _15473_/S vssd1 vssd1 vccd1 vccd1 _15468_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17206_ _25928_/Q _25994_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17207_/B sky130_fd_sc_hd__mux2_1
X_14418_ _14436_/A vssd1 vssd1 vccd1 vccd1 _14426_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_191_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18186_ _26279_/Q _26247_/Q _26215_/Q _26183_/Q _18185_/X _18068_/X vssd1 vssd1 vccd1
+ vccd1 _18186_/X sky130_fd_sc_hd__mux4_2
X_15398_ _15398_/A vssd1 vssd1 vccd1 vccd1 _26270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ _27076_/Q _27108_/Q _17173_/S vssd1 vssd1 vccd1 vccd1 _17137_/X sky130_fd_sc_hd__mux2_1
X_14349_ _26675_/Q _14337_/X _14345_/X _14348_/Y vssd1 vssd1 vccd1 vccd1 _26675_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17068_ _17068_/A vssd1 vssd1 vccd1 vccd1 _27920_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_144_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16019_ _16014_/Y _16015_/X _16016_/X _16017_/Y _16018_/X vssd1 vssd1 vccd1 vccd1
+ _16030_/C sky130_fd_sc_hd__a221o_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater400 _27266_/CLK vssd1 vssd1 vccd1 vccd1 _27576_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater411 _25958_/CLK vssd1 vssd1 vccd1 vccd1 _26051_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater422 _27327_/CLK vssd1 vssd1 vccd1 vccd1 _27323_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater433 _17407_/Y vssd1 vssd1 vccd1 vccd1 _26062_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19709_ _19709_/A vssd1 vssd1 vccd1 vccd1 _19709_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20981_ _20972_/X _20974_/X _20976_/X _20978_/X _20979_/X _20980_/X vssd1 vssd1 vccd1
+ vccd1 _20982_/A sky130_fd_sc_hd__mux4_1
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22720_ _22785_/A vssd1 vssd1 vccd1 vccd1 _22720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22651_ _22699_/A vssd1 vssd1 vccd1 vccd1 _22651_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21602_ _21650_/A vssd1 vssd1 vccd1 vccd1 _21602_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25370_ _25370_/A vssd1 vssd1 vccd1 vccd1 _27725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22582_ _22598_/A vssd1 vssd1 vccd1 vccd1 _22582_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24321_ _24321_/A vssd1 vssd1 vccd1 vccd1 _27444_/D sky130_fd_sc_hd__clkbuf_1
X_21533_ _21549_/A vssd1 vssd1 vccd1 vccd1 _21533_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27040_ _22946_/X _27040_/D vssd1 vssd1 vccd1 vccd1 _27040_/Q sky130_fd_sc_hd__dfxtp_1
X_24252_ _24330_/A vssd1 vssd1 vccd1 vccd1 _24287_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_21464_ _21464_/A vssd1 vssd1 vccd1 vccd1 _21464_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_153_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23203_ _23203_/A vssd1 vssd1 vccd1 vccd1 _27138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20415_ _20415_/A vssd1 vssd1 vccd1 vccd1 _20415_/X sky130_fd_sc_hd__clkbuf_1
X_21395_ _21653_/A vssd1 vssd1 vccd1 vccd1 _21464_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_24183_ _24183_/A vssd1 vssd1 vccd1 vccd1 _27362_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23134_ _23180_/S vssd1 vssd1 vccd1 vccd1 _23143_/S sky130_fd_sc_hd__clkbuf_2
X_20346_ _20334_/X _20335_/X _20336_/X _20337_/X _20339_/X _20341_/X vssd1 vssd1 vccd1
+ vccd1 _20347_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23065_ _23065_/A vssd1 vssd1 vccd1 vccd1 _27077_/D sky130_fd_sc_hd__clkbuf_1
X_20277_ _20277_/A vssd1 vssd1 vccd1 vccd1 _20277_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27942_ _27942_/A _15935_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_191_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22016_ _22083_/A vssd1 vssd1 vccd1 vccd1 _22016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26824_ _22192_/X _26824_/D vssd1 vssd1 vccd1 vccd1 _26824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26755_ _21956_/X _26755_/D vssd1 vssd1 vccd1 vccd1 _26755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23967_ _24014_/A vssd1 vssd1 vccd1 vccd1 _23967_/X sky130_fd_sc_hd__buf_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13720_ _26890_/Q _13710_/X _13718_/X _13719_/Y vssd1 vssd1 vccd1 vccd1 _26890_/D
+ sky130_fd_sc_hd__a31o_1
X_25706_ _25722_/A vssd1 vssd1 vccd1 vccd1 _25706_/X sky130_fd_sc_hd__clkbuf_1
X_22918_ _22918_/A vssd1 vssd1 vccd1 vccd1 _22918_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26686_ _21714_/X _26686_/D vssd1 vssd1 vccd1 vccd1 _26686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23898_ _27841_/Q _27145_/Q _25890_/Q _25858_/Q _23873_/X _23897_/X vssd1 vssd1 vccd1
+ vccd1 _23898_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13651_ _26914_/Q _13639_/X _13642_/X _13650_/Y vssd1 vssd1 vccd1 vccd1 _26914_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_95_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25637_ _25637_/A vssd1 vssd1 vccd1 vccd1 _25637_/X sky130_fd_sc_hd__clkbuf_1
X_22849_ _22837_/X _22838_/X _22839_/X _22840_/X _22841_/X _22842_/X vssd1 vssd1 vccd1
+ vccd1 _22850_/A sky130_fd_sc_hd__mux4_1
XFILLER_140_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16370_ _16359_/A _16357_/A _16369_/X vssd1 vssd1 vccd1 vccd1 _16371_/B sky130_fd_sc_hd__o21a_1
X_13582_ _14531_/A vssd1 vssd1 vccd1 vccd1 _13940_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25568_ _25568_/A vssd1 vssd1 vccd1 vccd1 _25568_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15321_/A vssd1 vssd1 vccd1 vccd1 _26304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27307_ _27308_/CLK _27307_/D vssd1 vssd1 vccd1 vccd1 _27307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24519_ _27608_/Q _24554_/B vssd1 vssd1 vccd1 vccd1 _24520_/A sky130_fd_sc_hd__and2_1
XFILLER_40_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25499_ _27700_/Q _25479_/X _25480_/X vssd1 vssd1 vccd1 vccd1 _25499_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_184_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _17972_/X _18033_/X _18039_/X _17932_/X vssd1 vssd1 vccd1 vccd1 _18052_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_40_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15252_ _14798_/X _26334_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15253_/A sky130_fd_sc_hd__mux2_1
X_27238_ _27258_/CLK _27238_/D vssd1 vssd1 vccd1 vccd1 _27238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ _14381_/A _14213_/B vssd1 vssd1 vccd1 vccd1 _14203_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15183_ _15183_/A vssd1 vssd1 vccd1 vccd1 _26365_/D sky130_fd_sc_hd__clkbuf_1
X_27169_ _27563_/CLK _27169_/D vssd1 vssd1 vccd1 vccd1 _27169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _14399_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14134_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19991_ _19991_/A vssd1 vssd1 vccd1 vccd1 _19991_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ _14079_/A vssd1 vssd1 vccd1 vccd1 _14070_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18942_ _18775_/X _18940_/X _18941_/X vssd1 vssd1 vccd1 vccd1 _18942_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13016_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13017_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18873_ _26684_/Q _26652_/Q _26620_/Q _26588_/Q _18847_/X _18782_/X vssd1 vssd1 vccd1
+ vccd1 _18873_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17824_ _17959_/A vssd1 vssd1 vccd1 vccd1 _17824_/X sky130_fd_sc_hd__buf_2
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17755_ _17755_/A vssd1 vssd1 vccd1 vccd1 _25936_/D sky130_fd_sc_hd__clkbuf_1
X_14967_ _26455_/Q _14957_/X _14960_/X _14966_/Y vssd1 vssd1 vccd1 vccd1 _26455_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16706_ _16619_/A _16703_/X _16705_/X vssd1 vssd1 vccd1 vccd1 _25618_/A sky130_fd_sc_hd__a21oi_2
X_13918_ _26819_/Q _13906_/X _13912_/X _13917_/Y vssd1 vssd1 vccd1 vccd1 _26819_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_130_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14898_ _14955_/S vssd1 vssd1 vccd1 vccd1 _14907_/S sky130_fd_sc_hd__clkbuf_2
X_17686_ _27411_/Q vssd1 vssd1 vccd1 vccd1 _17686_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19425_ _19419_/X _19421_/X _19424_/X _19290_/X _19360_/X vssd1 vssd1 vccd1 vccd1
+ _19426_/C sky130_fd_sc_hd__a221o_1
X_16637_ _16888_/A _16571_/X _16573_/X vssd1 vssd1 vccd1 vccd1 _16638_/B sky130_fd_sc_hd__a21o_1
X_13849_ _27270_/Q vssd1 vssd1 vccd1 vccd1 _15695_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19356_ _26415_/Q _26383_/Q _26351_/Q _26319_/Q _19331_/X _19240_/X vssd1 vssd1 vccd1
+ vccd1 _19356_/X sky130_fd_sc_hd__mux4_1
X_16568_ _16798_/B _16572_/B vssd1 vssd1 vccd1 vccd1 _16569_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18307_ _18304_/X _18306_/X _18331_/S vssd1 vssd1 vccd1 vccd1 _18307_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15519_ _13156_/X _26216_/Q _15523_/S vssd1 vssd1 vccd1 vccd1 _15520_/A sky130_fd_sc_hd__mux2_1
X_16499_ _16499_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16500_/B sky130_fd_sc_hd__and2_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19287_ _19287_/A vssd1 vssd1 vccd1 vccd1 _19287_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18238_ _18238_/A vssd1 vssd1 vccd1 vccd1 _18238_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1057 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18169_ _18161_/X _18164_/X _18167_/X _18168_/X _18122_/X vssd1 vssd1 vccd1 vccd1
+ _18170_/C sky130_fd_sc_hd__a221o_1
X_27994__460 vssd1 vssd1 vccd1 vccd1 _27994__460/HI _27994_/A sky130_fd_sc_hd__conb_1
XFILLER_7_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20200_ _20248_/A vssd1 vssd1 vccd1 vccd1 _20200_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21180_ _21212_/A vssd1 vssd1 vccd1 vccd1 _21180_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20131_ _20163_/A vssd1 vssd1 vccd1 vccd1 _20131_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_539 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20062_ _20078_/A vssd1 vssd1 vccd1 vccd1 _20062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24870_ _24889_/A _24870_/B vssd1 vssd1 vccd1 vccd1 _24870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_434 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater230 _26062_/CLK vssd1 vssd1 vccd1 vccd1 _26073_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater241 _27752_/CLK vssd1 vssd1 vccd1 vccd1 _27744_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater252 _27621_/CLK vssd1 vssd1 vccd1 vccd1 _27627_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23821_ _27072_/Q _27104_/Q _23845_/S vssd1 vssd1 vccd1 vccd1 _23821_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater263 _27172_/CLK vssd1 vssd1 vccd1 vccd1 _27607_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater274 _27372_/CLK vssd1 vssd1 vccd1 vccd1 _27475_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater285 _27480_/CLK vssd1 vssd1 vccd1 vccd1 _27484_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater296 _27263_/CLK vssd1 vssd1 vccd1 vccd1 _27245_/CLK sky130_fd_sc_hd__clkbuf_1
X_26540_ _21202_/X _26540_/D vssd1 vssd1 vccd1 vccd1 _26540_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 _18055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23752_ _24045_/S vssd1 vssd1 vccd1 vccd1 _23795_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 _18999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20964_ _20964_/A vssd1 vssd1 vccd1 vccd1 _20964_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22703_ _22961_/A vssd1 vssd1 vccd1 vccd1 _22772_/A sky130_fd_sc_hd__buf_2
X_26471_ _20964_/X _26471_/D vssd1 vssd1 vccd1 vccd1 _26471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23683_ _27767_/Q _27247_/Q _23683_/S vssd1 vssd1 vccd1 vccd1 _23684_/A sky130_fd_sc_hd__mux2_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ _20886_/X _20888_/X _20890_/X _20892_/X _20893_/X _20894_/X vssd1 vssd1 vccd1
+ vccd1 _20896_/A sky130_fd_sc_hd__mux4_1
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25422_ _27749_/Q input61/X _25424_/S vssd1 vssd1 vccd1 vccd1 _25423_/A sky130_fd_sc_hd__mux2_1
X_27962__448 vssd1 vssd1 vccd1 vccd1 _27962__448/HI _27962_/A sky130_fd_sc_hd__conb_1
X_22634_ _22699_/A vssd1 vssd1 vccd1 vccd1 _22634_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25353_ _25350_/A _25350_/B _25348_/A vssd1 vssd1 vccd1 vccd1 _25355_/A sky130_fd_sc_hd__o21ai_1
XFILLER_139_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22565_ _22597_/A vssd1 vssd1 vccd1 vccd1 _22565_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24304_ _24304_/A vssd1 vssd1 vccd1 vccd1 _24384_/B sky130_fd_sc_hd__clkbuf_4
X_21516_ _21564_/A vssd1 vssd1 vccd1 vccd1 _21516_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25284_ _27710_/Q _25263_/X _25283_/Y _25254_/X vssd1 vssd1 vccd1 vccd1 _27710_/D
+ sky130_fd_sc_hd__o211a_1
X_22496_ _22496_/A vssd1 vssd1 vccd1 vccd1 _22496_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_186_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27023_ _22884_/X _27023_/D vssd1 vssd1 vccd1 vccd1 _27023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24235_ _24235_/A _24235_/B vssd1 vssd1 vccd1 vccd1 _27389_/D sky130_fd_sc_hd__nor2_1
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21447_ _21463_/A vssd1 vssd1 vccd1 vccd1 _21447_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24166_ _24166_/A vssd1 vssd1 vccd1 vccd1 _27354_/D sky130_fd_sc_hd__clkbuf_1
X_21378_ _21378_/A vssd1 vssd1 vccd1 vccd1 _21378_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23117_ _27100_/Q _17683_/X _23121_/S vssd1 vssd1 vccd1 vccd1 _23118_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20329_ _20329_/A vssd1 vssd1 vccd1 vccd1 _20329_/X sky130_fd_sc_hd__clkbuf_1
X_24097_ _24119_/A vssd1 vssd1 vccd1 vccd1 _24106_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27925_ _27925_/A _15961_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
X_23048_ _27070_/Q _17689_/X _23048_/S vssd1 vssd1 vccd1 vccd1 _23049_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15870_ _15894_/A vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__buf_4
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27856_ _27856_/CLK _27856_/D vssd1 vssd1 vccd1 vccd1 _27856_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14821_ _14821_/A vssd1 vssd1 vccd1 vccd1 _26519_/D sky130_fd_sc_hd__clkbuf_1
X_26807_ _22136_/X _26807_/D vssd1 vssd1 vccd1 vccd1 _26807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27787_ _27787_/CLK _27787_/D vssd1 vssd1 vccd1 vccd1 _27787_/Q sky130_fd_sc_hd__dfxtp_1
X_24999_ _27965_/A _24998_/X _25024_/S vssd1 vssd1 vccd1 vccd1 _25000_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14752_ _14752_/A vssd1 vssd1 vccd1 vccd1 _26541_/D sky130_fd_sc_hd__clkbuf_1
X_17540_ _17437_/X _25847_/Q _17540_/S vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__mux2_1
X_26738_ _21892_/X _26738_/D vssd1 vssd1 vccd1 vccd1 _26738_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13884_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13703_/Y sky130_fd_sc_hd__nor2_1
X_17471_ _17471_/A vssd1 vssd1 vccd1 vccd1 _25825_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26669_ _21646_/X _26669_/D vssd1 vssd1 vccd1 vccd1 _26669_/Q sky130_fd_sc_hd__dfxtp_1
X_14683_ _26564_/Q _14671_/X _14679_/X _14682_/Y vssd1 vssd1 vccd1 vccd1 _26564_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_71_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19210_ _27808_/Q _26569_/Q _26441_/Q _26121_/Q _19118_/X _19183_/X vssd1 vssd1 vccd1
+ vccd1 _19210_/X sky130_fd_sc_hd__mux4_2
X_13634_ _13904_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13634_/Y sky130_fd_sc_hd__nor2_1
X_16422_ _16422_/A vssd1 vssd1 vccd1 vccd1 _16772_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19141_ _19299_/A vssd1 vssd1 vccd1 vccd1 _19261_/A sky130_fd_sc_hd__clkbuf_1
X_16353_ _16353_/A vssd1 vssd1 vccd1 vccd1 _16508_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_201_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13565_ _13930_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13565_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15304_ _26311_/Q _13379_/X _15306_/S vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__mux2_1
X_19072_ _19123_/A _19072_/B vssd1 vssd1 vccd1 vccd1 _19072_/X sky130_fd_sc_hd__or2_1
X_16284_ _16282_/Y _16119_/A _16277_/B _16536_/A _16283_/Y vssd1 vssd1 vccd1 vccd1
+ _24297_/A sky130_fd_sc_hd__o221a_1
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _27353_/Q _13062_/A _13082_/A _27321_/Q _13131_/X vssd1 vssd1 vccd1 vccd1
+ _16277_/A sky130_fd_sc_hd__a221oi_4
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15235_ _15235_/A vssd1 vssd1 vccd1 vccd1 _26342_/D sky130_fd_sc_hd__clkbuf_1
X_18023_ _26528_/Q _26496_/Q _26464_/Q _27040_/Q _17964_/X _17986_/X vssd1 vssd1 vccd1
+ vccd1 _18023_/X sky130_fd_sc_hd__mux4_1
X_15166_ _15166_/A vssd1 vssd1 vccd1 vccd1 _26373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ _14157_/A vssd1 vssd1 vccd1 vccd1 _14117_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15097_ _14782_/X _26403_/Q _15101_/S vssd1 vssd1 vccd1 vccd1 _15098_/A sky130_fd_sc_hd__mux2_1
X_19974_ _19990_/A vssd1 vssd1 vccd1 vccd1 _19974_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ _26782_/Q _14042_/X _14038_/X _14047_/Y vssd1 vssd1 vccd1 vccd1 _26782_/D
+ sky130_fd_sc_hd__a31o_1
X_18925_ _18921_/X _18924_/X _19553_/S vssd1 vssd1 vccd1 vccd1 _18925_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18856_ _19299_/A vssd1 vssd1 vccd1 vccd1 _19004_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_67_456 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17807_ _27593_/Q vssd1 vssd1 vccd1 vccd1 _18177_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_404 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18787_ _19297_/A vssd1 vssd1 vccd1 vccd1 _19208_/A sky130_fd_sc_hd__buf_2
X_15999_ _27482_/Q _27373_/Q vssd1 vssd1 vccd1 vccd1 _16001_/C sky130_fd_sc_hd__xnor2_1
X_17738_ _25931_/Q _17737_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17739_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17669_ _17520_/X _25905_/Q _17671_/S vssd1 vssd1 vccd1 vccd1 _17670_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19408_ _26834_/Q _26802_/Q _26770_/Q _26738_/Q _19338_/X _19407_/X vssd1 vssd1 vccd1
+ vccd1 _19409_/B sky130_fd_sc_hd__mux4_2
XFILLER_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20680_ _20668_/X _20669_/X _20670_/X _20671_/X _20672_/X _20673_/X vssd1 vssd1 vccd1
+ vccd1 _20681_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19339_ _26831_/Q _26799_/Q _26767_/Q _26735_/Q _19338_/X _19248_/X vssd1 vssd1 vccd1
+ vccd1 _19340_/B sky130_fd_sc_hd__mux4_2
XFILLER_148_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22350_ _22350_/A vssd1 vssd1 vccd1 vccd1 _22350_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21301_ _21301_/A vssd1 vssd1 vccd1 vccd1 _21301_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22281_ _22453_/A vssd1 vssd1 vccd1 vccd1 _22348_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24020_ _27093_/Q _24001_/X _24002_/X _27125_/Q _24003_/X vssd1 vssd1 vccd1 vccd1
+ _24020_/X sky130_fd_sc_hd__a221o_1
X_21232_ _22540_/A vssd1 vssd1 vccd1 vccd1 _21581_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21163_ _21211_/A vssd1 vssd1 vccd1 vccd1 _21163_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20114_ _20162_/A vssd1 vssd1 vccd1 vccd1 _20114_/X sky130_fd_sc_hd__clkbuf_1
X_25971_ _26068_/CLK _25971_/D vssd1 vssd1 vccd1 vccd1 _25971_/Q sky130_fd_sc_hd__dfxtp_1
X_21094_ _21126_/A vssd1 vssd1 vccd1 vccd1 _21094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27710_ _27770_/CLK _27710_/D vssd1 vssd1 vccd1 vccd1 _27710_/Q sky130_fd_sc_hd__dfxtp_1
X_20045_ _20077_/A vssd1 vssd1 vccd1 vccd1 _20045_/X sky130_fd_sc_hd__clkbuf_1
X_24922_ _24925_/B _24925_/C vssd1 vssd1 vccd1 vccd1 _24923_/B sky130_fd_sc_hd__xnor2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27641_ _27756_/CLK _27641_/D vssd1 vssd1 vccd1 vccd1 _27641_/Q sky130_fd_sc_hd__dfxtp_1
X_24853_ _24857_/B _24853_/B vssd1 vssd1 vccd1 vccd1 _24854_/B sky130_fd_sc_hd__or2_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23804_ _23946_/A vssd1 vssd1 vccd1 vccd1 _23804_/X sky130_fd_sc_hd__buf_2
XFILLER_2_1124 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27572_ _27572_/CLK _27572_/D vssd1 vssd1 vccd1 vccd1 _27572_/Q sky130_fd_sc_hd__dfxtp_1
X_24784_ _24841_/A vssd1 vssd1 vccd1 vccd1 _24861_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _19490_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21996_ _21996_/A vssd1 vssd1 vccd1 vccd1 _21996_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_116 _22540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _22616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26523_ _21140_/X _26523_/D vssd1 vssd1 vccd1 vccd1 _26523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _15773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23735_ _23735_/A vssd1 vssd1 vccd1 vccd1 _27269_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _20937_/X _20938_/X _20939_/X _20940_/X _20941_/X _20942_/X vssd1 vssd1 vccd1
+ vccd1 _20948_/A sky130_fd_sc_hd__mux4_1
XANTENNA_149 _13133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26454_ _20904_/X _26454_/D vssd1 vssd1 vccd1 vccd1 _26454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23666_ _24848_/A _27239_/Q _23672_/S vssd1 vssd1 vccd1 vccd1 _23667_/A sky130_fd_sc_hd__mux2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20878_ _20878_/A vssd1 vssd1 vccd1 vccd1 _20878_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25405_ _27741_/Q input53/X _25413_/S vssd1 vssd1 vccd1 vccd1 _25406_/A sky130_fd_sc_hd__mux2_1
X_22617_ _22961_/A vssd1 vssd1 vccd1 vccd1 _22686_/A sky130_fd_sc_hd__buf_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26385_ _20659_/X _26385_/D vssd1 vssd1 vccd1 vccd1 _26385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23597_ _23597_/A vssd1 vssd1 vccd1 vccd1 _27219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25336_ _25344_/A _25336_/B vssd1 vssd1 vccd1 vccd1 _25336_/Y sky130_fd_sc_hd__nand2_1
X_13350_ _14740_/A vssd1 vssd1 vccd1 vccd1 _13350_/X sky130_fd_sc_hd__clkbuf_4
X_22548_ _22612_/A vssd1 vssd1 vccd1 vccd1 _22548_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25267_ _25267_/A _25267_/B vssd1 vssd1 vccd1 vccd1 _25267_/Y sky130_fd_sc_hd__nor2_1
X_13281_ _13281_/A vssd1 vssd1 vccd1 vccd1 _27019_/D sky130_fd_sc_hd__clkbuf_1
X_22479_ _22471_/X _22472_/X _22473_/X _22474_/X _22475_/X _22476_/X vssd1 vssd1 vccd1
+ vccd1 _22480_/A sky130_fd_sc_hd__mux4_1
X_15020_ _26436_/Q _15015_/X _15016_/X _15019_/Y vssd1 vssd1 vccd1 vccd1 _26436_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27006_ _22830_/X _27006_/D vssd1 vssd1 vccd1 vccd1 _27006_/Q sky130_fd_sc_hd__dfxtp_1
X_24218_ _24218_/A _24222_/B vssd1 vssd1 vccd1 vccd1 _27377_/D sky130_fd_sc_hd__nor2_1
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25198_ _25198_/A _25198_/B vssd1 vssd1 vccd1 vccd1 _25199_/B sky130_fd_sc_hd__xor2_1
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24149_ _27452_/Q _24151_/B vssd1 vssd1 vccd1 vccd1 _24150_/A sky130_fd_sc_hd__and2_1
XFILLER_122_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16971_ _16979_/B _16971_/B vssd1 vssd1 vccd1 vccd1 _16982_/D sky130_fd_sc_hd__and2_1
XFILLER_7_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18710_ _18710_/A vssd1 vssd1 vccd1 vccd1 _26017_/D sky130_fd_sc_hd__clkbuf_1
X_15922_ _15924_/A vssd1 vssd1 vccd1 vccd1 _15922_/Y sky130_fd_sc_hd__inv_2
X_19690_ _19678_/X _19679_/X _19680_/X _19681_/X _19682_/X _19683_/X vssd1 vssd1 vccd1
+ vccd1 _19691_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18641_ _25987_/Q _17705_/X _18641_/S vssd1 vssd1 vccd1 vccd1 _18642_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27839_ _27840_/CLK _27839_/D vssd1 vssd1 vccd1 vccd1 _27839_/Q sky130_fd_sc_hd__dfxtp_1
X_15853_ _13240_/X _26074_/Q _15853_/S vssd1 vssd1 vccd1 vccd1 _15854_/A sky130_fd_sc_hd__mux2_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14804_ _14804_/A vssd1 vssd1 vccd1 vccd1 _14804_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _18009_/X _18569_/X _18571_/X _18014_/X vssd1 vssd1 vccd1 vccd1 _18572_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _27800_/Q _12998_/B vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__and2_1
XFILLER_18_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15784_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15853_/S sky130_fd_sc_hd__buf_2
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _27439_/Q vssd1 vssd1 vccd1 vccd1 _17523_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14735_ _14734_/X _26546_/Q _14741_/S vssd1 vssd1 vccd1 vccd1 _14736_/A sky130_fd_sc_hd__mux2_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14666_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _17453_/X _25820_/Q _17454_/S vssd1 vssd1 vccd1 vccd1 _17455_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13617_ _13887_/A _13621_/B vssd1 vssd1 vccd1 vccd1 _13617_/Y sky130_fd_sc_hd__nor2_1
X_16405_ _16774_/B vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14597_ _15758_/A _14597_/B vssd1 vssd1 vccd1 vccd1 _14597_/Y sky130_fd_sc_hd__nor2_1
X_17385_ _27097_/Q _27129_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17385_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19124_ _26277_/Q _26245_/Q _26213_/Q _26181_/Q _19028_/X _19074_/X vssd1 vssd1 vccd1
+ vccd1 _19124_/X sky130_fd_sc_hd__mux4_2
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13548_ _26946_/Q _13535_/X _13528_/X _13547_/Y vssd1 vssd1 vccd1 vccd1 _26946_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_146_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16336_ _16756_/A _16336_/B vssd1 vssd1 vccd1 vccd1 _16349_/B sky130_fd_sc_hd__xnor2_1
XFILLER_146_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ _16266_/A _24293_/A _16266_/Y vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__o21ai_1
X_19055_ _26402_/Q _26370_/Q _26338_/Q _26306_/Q _19054_/X _18982_/X vssd1 vssd1 vccd1
+ vccd1 _19055_/X sky130_fd_sc_hd__mux4_1
X_13479_ _14452_/A vssd1 vssd1 vccd1 vccd1 _13884_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18006_ _26688_/Q _26656_/Q _26624_/Q _26592_/Q _18004_/X _18005_/X vssd1 vssd1 vccd1
+ vccd1 _18008_/A sky130_fd_sc_hd__mux4_2
X_15218_ _15218_/A vssd1 vssd1 vccd1 vccd1 _26350_/D sky130_fd_sc_hd__clkbuf_1
X_16198_ _27522_/Q _15991_/A vssd1 vssd1 vccd1 vccd1 _16198_/X sky130_fd_sc_hd__or2b_1
XFILLER_126_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ _26380_/Q _13363_/X _15151_/S vssd1 vssd1 vccd1 vccd1 _15150_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19957_ _19989_/A vssd1 vssd1 vccd1 vccd1 _19957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18908_ _19441_/A vssd1 vssd1 vccd1 vccd1 _18908_/X sky130_fd_sc_hd__buf_4
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19888_ _19882_/X _19883_/X _19884_/X _19885_/X _19886_/X _19887_/X vssd1 vssd1 vccd1
+ vccd1 _19889_/A sky130_fd_sc_hd__mux4_1
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18839_ _19469_/A vssd1 vssd1 vccd1 vccd1 _19220_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21850_ _21914_/A vssd1 vssd1 vccd1 vccd1 _21850_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20801_ _22546_/A vssd1 vssd1 vccd1 vccd1 _21149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21781_ _21813_/A vssd1 vssd1 vccd1 vccd1 _21781_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23520_ _27756_/Q vssd1 vssd1 vccd1 vccd1 _24835_/B sky130_fd_sc_hd__buf_2
XFILLER_196_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20732_ _20722_/X _20723_/X _20724_/X _20725_/X _20726_/X _20727_/X vssd1 vssd1 vccd1
+ vccd1 _20733_/A sky130_fd_sc_hd__mux4_1
XFILLER_168_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23451_ _27174_/Q _23456_/B vssd1 vssd1 vccd1 vccd1 _23451_/X sky130_fd_sc_hd__or2_1
XFILLER_149_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20663_ _20663_/A vssd1 vssd1 vccd1 vccd1 _20663_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22402_ _22434_/A vssd1 vssd1 vccd1 vccd1 _22402_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26170_ _19907_/X _26170_/D vssd1 vssd1 vccd1 vccd1 _26170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23382_ _27762_/Q vssd1 vssd1 vccd1 vccd1 _24862_/A sky130_fd_sc_hd__buf_2
XFILLER_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20594_ _20582_/X _20583_/X _20584_/X _20585_/X _20586_/X _20587_/X vssd1 vssd1 vccd1
+ vccd1 _20595_/A sky130_fd_sc_hd__mux4_2
X_25121_ _25119_/X _25129_/A vssd1 vssd1 vccd1 vccd1 _25122_/B sky130_fd_sc_hd__and2b_1
X_22333_ _22349_/A vssd1 vssd1 vccd1 vccd1 _22333_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_567 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25052_ _27229_/Q vssd1 vssd1 vccd1 vccd1 _25052_/X sky130_fd_sc_hd__buf_2
X_22264_ _22264_/A vssd1 vssd1 vccd1 vccd1 _22264_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24003_ _24003_/A vssd1 vssd1 vccd1 vccd1 _24003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21215_ _21215_/A vssd1 vssd1 vccd1 vccd1 _21289_/A sky130_fd_sc_hd__buf_2
XFILLER_105_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22195_ _22453_/A vssd1 vssd1 vccd1 vccd1 _22262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21146_ _21212_/A vssd1 vssd1 vccd1 vccd1 _21146_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21077_ _21125_/A vssd1 vssd1 vccd1 vccd1 _21077_/X sky130_fd_sc_hd__clkbuf_1
X_25954_ _25958_/CLK _25954_/D vssd1 vssd1 vccd1 vccd1 _25954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24905_ _27657_/Q _24885_/X _24904_/Y _24890_/X vssd1 vssd1 vccd1 vccd1 _27657_/D
+ sky130_fd_sc_hd__o211a_1
X_20028_ _20076_/A vssd1 vssd1 vccd1 vccd1 _20028_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25885_ _25923_/CLK _25885_/D vssd1 vssd1 vccd1 vccd1 _25885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27624_ _27627_/CLK _27624_/D vssd1 vssd1 vccd1 vccd1 _27624_/Q sky130_fd_sc_hd__dfxtp_1
X_24836_ _24835_/B _24831_/B _24835_/A vssd1 vssd1 vccd1 vccd1 _24837_/B sky130_fd_sc_hd__a21oi_1
XFILLER_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24767_ _24767_/A _24772_/B vssd1 vssd1 vccd1 vccd1 _24767_/Y sky130_fd_sc_hd__nand2_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27555_ _27555_/CLK _27555_/D vssd1 vssd1 vccd1 vccd1 _27555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _21965_/X _21966_/X _21967_/X _21968_/X _21969_/X _21970_/X vssd1 vssd1 vccd1
+ vccd1 _21980_/A sky130_fd_sc_hd__mux4_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _26622_/Q _14514_/X _14510_/X _14519_/Y vssd1 vssd1 vccd1 vccd1 _26622_/D
+ sky130_fd_sc_hd__a31o_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23718_ _24965_/A _27263_/Q _23720_/S vssd1 vssd1 vccd1 vccd1 _23719_/A sky130_fd_sc_hd__mux2_1
X_26506_ _21086_/X _26506_/D vssd1 vssd1 vccd1 vccd1 _26506_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27486_ _27600_/CLK _27486_/D vssd1 vssd1 vccd1 vccd1 _27486_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24698_ _27181_/Q _24698_/B vssd1 vssd1 vccd1 vccd1 _24698_/X sky130_fd_sc_hd__or2_1
XFILLER_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _26641_/Q _14441_/X _14437_/X _14450_/Y vssd1 vssd1 vccd1 vccd1 _26641_/D
+ sky130_fd_sc_hd__a31o_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26437_ _20843_/X _26437_/D vssd1 vssd1 vccd1 vccd1 _26437_/Q sky130_fd_sc_hd__dfxtp_1
X_23649_ _23649_/A _23649_/B vssd1 vssd1 vccd1 vccd1 _27232_/D sky130_fd_sc_hd__nor2_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13402_ _13402_/A vssd1 vssd1 vccd1 vccd1 _13415_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17170_ _25824_/Q _26023_/Q _17219_/S vssd1 vssd1 vccd1 vccd1 _17170_/X sky130_fd_sc_hd__mux2_1
X_14382_ _26663_/Q _14379_/X _14371_/X _14381_/Y vssd1 vssd1 vccd1 vccd1 _26663_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26368_ _20595_/X _26368_/D vssd1 vssd1 vccd1 vccd1 _26368_/Q sky130_fd_sc_hd__dfxtp_1
X_16121_ _16277_/B vssd1 vssd1 vccd1 vccd1 _16121_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25319_ _25328_/A _25319_/B _25319_/C vssd1 vssd1 vccd1 vccd1 _25320_/B sky130_fd_sc_hd__and3_1
X_13333_ _13333_/A vssd1 vssd1 vccd1 vccd1 _26998_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26299_ _20351_/X _26299_/D vssd1 vssd1 vccd1 vccd1 _26299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16052_ _27477_/Q vssd1 vssd1 vccd1 vccd1 _16052_/Y sky130_fd_sc_hd__inv_2
X_13264_ _13264_/A vssd1 vssd1 vccd1 vccd1 _27027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15003_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15003_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13195_ _13231_/B vssd1 vssd1 vccd1 vccd1 _13237_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19811_ _19811_/A vssd1 vssd1 vccd1 vccd1 _19811_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19742_ _19726_/X _19727_/X _19728_/X _19729_/X _19731_/X _19733_/X vssd1 vssd1 vccd1
+ vccd1 _19743_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16954_ _27582_/Q vssd1 vssd1 vccd1 vccd1 _24635_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15905_ _15906_/A vssd1 vssd1 vccd1 vccd1 _15905_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19673_ _19673_/A vssd1 vssd1 vccd1 vccd1 _19673_/X sky130_fd_sc_hd__clkbuf_1
X_16885_ _16885_/A _16885_/B vssd1 vssd1 vccd1 vccd1 _16885_/X sky130_fd_sc_hd__xor2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18624_ _25979_/Q _17680_/X _18630_/S vssd1 vssd1 vccd1 vccd1 _18625_/A sky130_fd_sc_hd__mux2_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _13190_/X _26082_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15837_/A sky130_fd_sc_hd__mux2_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18555_ _18468_/X _18550_/X _18554_/X _18016_/X vssd1 vssd1 vccd1 vccd1 _18564_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _15767_/A _15771_/B vssd1 vssd1 vccd1 vccd1 _15767_/Y sky130_fd_sc_hd__nor2_1
X_12979_ _27808_/Q _12987_/B vssd1 vssd1 vccd1 vccd1 _12980_/A sky130_fd_sc_hd__and2_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17506_ _17504_/X _25836_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17507_/A sky130_fd_sc_hd__mux2_1
X_14718_ _14718_/A vssd1 vssd1 vccd1 vccd1 _14718_/X sky130_fd_sc_hd__buf_2
XFILLER_162_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18486_ _18486_/A vssd1 vssd1 vccd1 vccd1 _18486_/X sky130_fd_sc_hd__clkbuf_2
X_15698_ _15712_/A vssd1 vssd1 vccd1 vccd1 _15703_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17437_ _27412_/Q vssd1 vssd1 vccd1 vccd1 _17437_/X sky130_fd_sc_hd__clkbuf_1
X_14649_ _15723_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14649_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_16 _25992_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_27 _27143_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 _18481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17368_ _17368_/A vssd1 vssd1 vccd1 vccd1 _27945_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19107_ _19107_/A _19107_/B _19107_/C vssd1 vssd1 vccd1 vccd1 _19108_/A sky130_fd_sc_hd__and3_1
X_16319_ _16836_/A _16319_/B vssd1 vssd1 vccd1 vccd1 _16598_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17299_ _17299_/A vssd1 vssd1 vccd1 vccd1 _17299_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19038_ _19038_/A vssd1 vssd1 vccd1 vccd1 _26049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21000_ _21000_/A vssd1 vssd1 vccd1 vccd1 _21000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22951_ _22939_/X _22940_/X _22941_/X _22942_/X _22943_/X _22944_/X vssd1 vssd1 vccd1
+ vccd1 _22952_/A sky130_fd_sc_hd__mux4_1
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21902_ _21902_/A vssd1 vssd1 vccd1 vccd1 _21902_/X sky130_fd_sc_hd__clkbuf_1
X_25670_ _25670_/A vssd1 vssd1 vccd1 vccd1 _25670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22882_ _22882_/A vssd1 vssd1 vccd1 vccd1 _22882_/X sky130_fd_sc_hd__clkbuf_1
X_24621_ _24621_/A vssd1 vssd1 vccd1 vccd1 _27569_/D sky130_fd_sc_hd__clkbuf_1
X_21833_ _21825_/X _21826_/X _21827_/X _21828_/X _21830_/X _21832_/X vssd1 vssd1 vccd1
+ vccd1 _21834_/A sky130_fd_sc_hd__mux4_1
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27340_ _27342_/CLK _27340_/D vssd1 vssd1 vccd1 vccd1 _27340_/Q sky130_fd_sc_hd__dfxtp_2
X_24552_ _24552_/A _24552_/B vssd1 vssd1 vccd1 vccd1 _24553_/A sky130_fd_sc_hd__and2_1
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21764_ _21828_/A vssd1 vssd1 vccd1 vccd1 _21764_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23503_ _27194_/Q _23650_/B vssd1 vssd1 vccd1 vccd1 _23503_/X sky130_fd_sc_hd__or2_1
XFILLER_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20715_ _20715_/A vssd1 vssd1 vccd1 vccd1 _20715_/X sky130_fd_sc_hd__clkbuf_1
X_27271_ _27410_/CLK _27271_/D vssd1 vssd1 vccd1 vccd1 _27271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24483_ _27638_/Q _24509_/B vssd1 vssd1 vccd1 vccd1 _24484_/A sky130_fd_sc_hd__and2_1
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21695_ _21689_/X _21690_/X _21691_/X _21692_/X _21693_/X _21694_/X vssd1 vssd1 vccd1
+ vccd1 _21696_/A sky130_fd_sc_hd__mux4_1
X_26222_ _20089_/X _26222_/D vssd1 vssd1 vccd1 vccd1 _26222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23434_ _23624_/A vssd1 vssd1 vccd1 vccd1 _23434_/X sky130_fd_sc_hd__clkbuf_2
X_20646_ _20636_/X _20637_/X _20638_/X _20639_/X _20640_/X _20641_/X vssd1 vssd1 vccd1
+ vccd1 _20647_/A sky130_fd_sc_hd__mux4_1
X_26153_ _19847_/X _26153_/D vssd1 vssd1 vccd1 vccd1 _26153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23365_ _27251_/Q vssd1 vssd1 vccd1 vccd1 _23365_/Y sky130_fd_sc_hd__inv_2
X_20577_ _20577_/A vssd1 vssd1 vccd1 vccd1 _20577_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25104_ _27978_/A _25103_/X _25104_/S vssd1 vssd1 vccd1 vccd1 _25105_/A sky130_fd_sc_hd__mux2_1
XFILLER_178_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22316_ _22348_/A vssd1 vssd1 vccd1 vccd1 _22316_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26084_ _19604_/X _26084_/D vssd1 vssd1 vccd1 vccd1 _26084_/Q sky130_fd_sc_hd__dfxtp_1
X_23296_ input46/X vssd1 vssd1 vccd1 vccd1 _23296_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25035_ _25035_/A vssd1 vssd1 vccd1 vccd1 _25035_/X sky130_fd_sc_hd__clkbuf_2
X_22247_ _22263_/A vssd1 vssd1 vccd1 vccd1 _22247_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22178_ _22523_/A vssd1 vssd1 vccd1 vccd1 _22249_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21129_ _21215_/A vssd1 vssd1 vccd1 vccd1 _21199_/A sky130_fd_sc_hd__buf_2
X_26986_ _22760_/X _26986_/D vssd1 vssd1 vccd1 vccd1 _26986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25937_ _27851_/CLK _25937_/D vssd1 vssd1 vccd1 vccd1 _25937_/Q sky130_fd_sc_hd__dfxtp_1
X_13951_ _14333_/A _13954_/B vssd1 vssd1 vccd1 vccd1 _13951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13882_ _13882_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13882_/Y sky130_fd_sc_hd__nor2_1
X_16670_ _16670_/A _16809_/B vssd1 vssd1 vccd1 vccd1 _16670_/Y sky130_fd_sc_hd__nor2_1
X_25868_ _25901_/CLK _25868_/D vssd1 vssd1 vccd1 vccd1 _25868_/Q sky130_fd_sc_hd__dfxtp_1
X_27607_ _27607_/CLK _27607_/D vssd1 vssd1 vccd1 vccd1 _27607_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _26170_/Q _14810_/A _15621_/S vssd1 vssd1 vccd1 vccd1 _15622_/A sky130_fd_sc_hd__mux2_1
X_24819_ _27784_/Q vssd1 vssd1 vccd1 vccd1 _24969_/A sky130_fd_sc_hd__inv_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25799_ _17514_/X _27854_/Q _25801_/S vssd1 vssd1 vccd1 vccd1 _25800_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _26958_/Q _26926_/Q _26894_/Q _26862_/Q _18011_/A _18427_/A vssd1 vssd1 vccd1
+ vccd1 _18340_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27538_ _27610_/CLK _27538_/D vssd1 vssd1 vccd1 vccd1 _27538_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15608_/A vssd1 vssd1 vccd1 vccd1 _15621_/S sky130_fd_sc_hd__buf_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14503_/A vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__clkbuf_2
X_18271_ _18268_/X _18270_/X _18378_/S vssd1 vssd1 vccd1 vccd1 _18271_/X sky130_fd_sc_hd__mux2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _15483_/A vssd1 vssd1 vccd1 vccd1 _26233_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27469_ _27472_/CLK _27469_/D vssd1 vssd1 vccd1 vccd1 _27469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17222_ _17177_/X _17215_/X _17218_/X _17221_/X vssd1 vssd1 vccd1 vccd1 _17222_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14434_ _15710_/A _14446_/B vssd1 vssd1 vccd1 vccd1 _14434_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_28003__469 vssd1 vssd1 vccd1 vccd1 _28003__469/HI _28003_/A sky130_fd_sc_hd__conb_1
Xinput14 la1_data_in[14] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14365_ _14365_/A vssd1 vssd1 vccd1 vccd1 _14365_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17153_ _17153_/A vssd1 vssd1 vccd1 vccd1 _27927_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 la1_data_in[24] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_2
Xinput36 la1_data_in[5] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput47 la1_oenb[15] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_4
Xinput58 la1_oenb[25] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_8
XFILLER_183_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13316_ _13316_/A vssd1 vssd1 vccd1 vccd1 _27003_/D sky130_fd_sc_hd__clkbuf_1
X_16104_ _16360_/A vssd1 vssd1 vccd1 vccd1 _16486_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 la1_oenb[6] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_6
XFILLER_155_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17084_ _25918_/Q _25984_/Q _17132_/S vssd1 vssd1 vccd1 vccd1 _17085_/B sky130_fd_sc_hd__mux2_1
X_14296_ _14296_/A vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13247_ _15783_/A _14813_/B vssd1 vssd1 vccd1 vccd1 _13304_/A sky130_fd_sc_hd__nor2_2
X_16035_ _16254_/S vssd1 vssd1 vccd1 vccd1 _16266_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13178_ _16169_/A vssd1 vssd1 vccd1 vccd1 _14779_/A sky130_fd_sc_hd__buf_2
XFILLER_112_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_401 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17986_ _18141_/A vssd1 vssd1 vccd1 vccd1 _17986_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19725_ _19725_/A vssd1 vssd1 vccd1 vccd1 _19725_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16937_ _27598_/Q vssd1 vssd1 vccd1 vccd1 _18828_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19656_ _19637_/X _19638_/X _19639_/X _19640_/X _19644_/X _19647_/X vssd1 vssd1 vccd1
+ vccd1 _19657_/A sky130_fd_sc_hd__mux4_1
X_16868_ _25909_/Q _16755_/A _16753_/B _16646_/B vssd1 vssd1 vccd1 vccd1 _16868_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18607_ _25976_/Q vssd1 vssd1 vccd1 vccd1 _24823_/A sky130_fd_sc_hd__inv_2
XFILLER_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15819_ _13144_/X _26090_/Q _15827_/S vssd1 vssd1 vccd1 vccd1 _15820_/A sky130_fd_sc_hd__mux2_1
X_19587_ _19570_/X _19572_/X _19574_/X _19576_/X _19577_/X _19578_/X vssd1 vssd1 vccd1
+ vccd1 _19588_/A sky130_fd_sc_hd__mux4_1
X_16799_ _16648_/X _16650_/B _16797_/X _16798_/Y vssd1 vssd1 vccd1 vccd1 _16800_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18538_ _26167_/Q _26103_/Q _27031_/Q _26999_/Q _18455_/X _18011_/X vssd1 vssd1 vccd1
+ vccd1 _18539_/A sky130_fd_sc_hd__mux4_2
X_18469_ _27819_/Q _26580_/Q _26452_/Q _26132_/Q _18401_/X _18425_/X vssd1 vssd1 vccd1
+ vccd1 _18469_/X sky130_fd_sc_hd__mux4_1
XFILLER_178_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20500_ _20500_/A vssd1 vssd1 vccd1 vccd1 _20500_/X sky130_fd_sc_hd__clkbuf_2
X_21480_ _21549_/A vssd1 vssd1 vccd1 vccd1 _21480_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20431_ _25641_/A vssd1 vssd1 vccd1 vccd1 _20776_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23150_ _27115_/Q _17731_/X _23154_/S vssd1 vssd1 vccd1 vccd1 _23151_/A sky130_fd_sc_hd__mux2_1
X_20362_ _20708_/A vssd1 vssd1 vccd1 vccd1 _20427_/A sky130_fd_sc_hd__buf_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22101_ _22537_/A vssd1 vssd1 vccd1 vccd1 _22451_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23081_ _27085_/Q _17737_/X _23081_/S vssd1 vssd1 vccd1 vccd1 _23082_/A sky130_fd_sc_hd__mux2_1
X_20293_ _20293_/A vssd1 vssd1 vccd1 vccd1 _20293_/X sky130_fd_sc_hd__clkbuf_1
X_22032_ _22032_/A vssd1 vssd1 vccd1 vccd1 _22032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_624 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26840_ _22252_/X _26840_/D vssd1 vssd1 vccd1 vccd1 _26840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23983_ _27850_/Q _27154_/Q _25899_/Q _25867_/Q _23967_/X _23944_/X vssd1 vssd1 vccd1
+ vccd1 _23983_/X sky130_fd_sc_hd__mux4_1
X_26771_ _22008_/X _26771_/D vssd1 vssd1 vccd1 vccd1 _26771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22934_ _22934_/A vssd1 vssd1 vccd1 vccd1 _22934_/X sky130_fd_sc_hd__clkbuf_1
X_25722_ _25722_/A vssd1 vssd1 vccd1 vccd1 _25722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25653_ _25653_/A vssd1 vssd1 vccd1 vccd1 _25721_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22865_ _22853_/X _22854_/X _22855_/X _22856_/X _22857_/X _22858_/X vssd1 vssd1 vccd1
+ vccd1 _22866_/A sky130_fd_sc_hd__mux4_1
XFILLER_189_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21816_ _21816_/A vssd1 vssd1 vccd1 vccd1 _21816_/X sky130_fd_sc_hd__clkbuf_1
X_24604_ _24604_/A vssd1 vssd1 vccd1 vccd1 _27561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25584_ _25584_/A vssd1 vssd1 vccd1 vccd1 _25584_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22796_ _22796_/A vssd1 vssd1 vccd1 vccd1 _22796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24535_ _24534_/X _16979_/A _24545_/S vssd1 vssd1 vccd1 vccd1 _24536_/B sky130_fd_sc_hd__mux2_1
X_27323_ _27323_/CLK _27323_/D vssd1 vssd1 vccd1 vccd1 _27323_/Q sky130_fd_sc_hd__dfxtp_1
X_21747_ _21737_/X _21738_/X _21739_/X _21740_/X _21743_/X _21746_/X vssd1 vssd1 vccd1
+ vccd1 _21748_/A sky130_fd_sc_hd__mux4_1
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27254_ _27781_/CLK _27254_/D vssd1 vssd1 vccd1 vccd1 _27254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24466_ _24466_/A vssd1 vssd1 vccd1 vccd1 _27509_/D sky130_fd_sc_hd__clkbuf_1
X_21678_ _21726_/A vssd1 vssd1 vccd1 vccd1 _21678_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_769 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23417_ _23485_/A vssd1 vssd1 vccd1 vccd1 _23500_/B sky130_fd_sc_hd__clkbuf_2
X_26205_ _20035_/X _26205_/D vssd1 vssd1 vccd1 vccd1 _26205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20629_ _20629_/A vssd1 vssd1 vccd1 vccd1 _20629_/X sky130_fd_sc_hd__clkbuf_1
X_27185_ _27185_/CLK _27185_/D vssd1 vssd1 vccd1 vccd1 _27185_/Q sky130_fd_sc_hd__dfxtp_1
X_24397_ _24397_/A vssd1 vssd1 vccd1 vccd1 _27478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14150_ _14166_/A vssd1 vssd1 vccd1 vccd1 _14234_/B sky130_fd_sc_hd__clkbuf_2
X_26136_ _19789_/X _26136_/D vssd1 vssd1 vccd1 vccd1 _26136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23348_ _27761_/Q vssd1 vssd1 vccd1 vccd1 _24754_/A sky130_fd_sc_hd__inv_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _13101_/A vssd1 vssd1 vccd1 vccd1 _27058_/D sky130_fd_sc_hd__clkbuf_1
X_14081_ _14346_/A _14085_/B vssd1 vssd1 vccd1 vccd1 _14081_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26067_ _26067_/CLK _26067_/D vssd1 vssd1 vccd1 vccd1 _26067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23279_ _23266_/Y input55/X _23276_/Y input56/X _23278_/X vssd1 vssd1 vccd1 vccd1
+ _23321_/A sky130_fd_sc_hd__a221o_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25018_ _25018_/A vssd1 vssd1 vccd1 vccd1 _25018_/X sky130_fd_sc_hd__buf_2
X_13032_ _13231_/B vssd1 vssd1 vccd1 vccd1 _13201_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17840_ _17898_/A vssd1 vssd1 vccd1 vccd1 _18392_/A sky130_fd_sc_hd__buf_2
XFILLER_105_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17771_ _17771_/A vssd1 vssd1 vccd1 vccd1 _25941_/D sky130_fd_sc_hd__clkbuf_1
X_14983_ _15023_/A vssd1 vssd1 vccd1 vccd1 _14994_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_26969_ _22696_/X _26969_/D vssd1 vssd1 vccd1 vccd1 _26969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19510_ _26550_/Q _26518_/Q _26486_/Q _27062_/Q _18896_/X _19445_/X vssd1 vssd1 vccd1
+ vccd1 _19510_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16722_ _16722_/A _16786_/B vssd1 vssd1 vccd1 vccd1 _16722_/X sky130_fd_sc_hd__or2_1
X_13934_ _13934_/A _13940_/B vssd1 vssd1 vccd1 vccd1 _13934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19441_ _19441_/A vssd1 vssd1 vccd1 vccd1 _19441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _16888_/A _16888_/B _16572_/X vssd1 vssd1 vccd1 vccd1 _16654_/B sky130_fd_sc_hd__a21o_1
X_13865_ _13919_/A vssd1 vssd1 vccd1 vccd1 _13865_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15604_ _26178_/Q _14785_/A _15606_/S vssd1 vssd1 vccd1 vccd1 _15605_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19372_ _18895_/X _19367_/X _19369_/X _19371_/X _19258_/X vssd1 vssd1 vccd1 vccd1
+ _19381_/B sky130_fd_sc_hd__a221o_1
X_16584_ _16831_/B _16588_/B vssd1 vssd1 vccd1 vccd1 _16584_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13796_ _26863_/Q _13793_/X _13794_/X _13795_/Y vssd1 vssd1 vccd1 vccd1 _26863_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_31_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18323_ _18323_/A _18322_/X vssd1 vssd1 vccd1 vccd1 _18323_/X sky130_fd_sc_hd__or2b_1
XFILLER_187_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15535_ _15535_/A vssd1 vssd1 vccd1 vccd1 _26209_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18254_ _18150_/X _18247_/X _18252_/X _18253_/X vssd1 vssd1 vccd1 vccd1 _18264_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15466_ _15466_/A vssd1 vssd1 vccd1 vccd1 _26240_/D sky130_fd_sc_hd__clkbuf_1
X_17205_ _17266_/A vssd1 vssd1 vccd1 vccd1 _17254_/S sky130_fd_sc_hd__clkbuf_2
X_14417_ _16033_/A vssd1 vssd1 vccd1 vccd1 _15699_/A sky130_fd_sc_hd__buf_2
XFILLER_8_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18185_ _18458_/A vssd1 vssd1 vccd1 vccd1 _18185_/X sky130_fd_sc_hd__buf_2
X_15397_ _14798_/X _26270_/Q _15401_/S vssd1 vssd1 vccd1 vccd1 _15398_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1037 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17136_ _17116_/X _17131_/X _17133_/X _17135_/X vssd1 vssd1 vccd1 vccd1 _17136_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14348_ _14348_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _14348_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14279_ _14367_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17067_ _27199_/Q _17066_/X _17067_/S vssd1 vssd1 vccd1 vccd1 _17068_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16018_ _27479_/Q _27266_/Q vssd1 vssd1 vccd1 vccd1 _16018_/X sky130_fd_sc_hd__xor2_1
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater401 _27338_/CLK vssd1 vssd1 vccd1 vccd1 _27266_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater412 _27386_/CLK vssd1 vssd1 vccd1 vccd1 _27388_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_100_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17969_ _17961_/X _17963_/X _17968_/X _17854_/X _17856_/X vssd1 vssd1 vccd1 vccd1
+ _17970_/C sky130_fd_sc_hd__a221o_1
XFILLER_100_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater423 _27328_/CLK vssd1 vssd1 vccd1 vccd1 _27327_/CLK sky130_fd_sc_hd__clkbuf_1
X_19708_ _19694_/X _19695_/X _19696_/X _19697_/X _19698_/X _19699_/X vssd1 vssd1 vccd1
+ vccd1 _19709_/A sky130_fd_sc_hd__mux4_1
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20980_ _21028_/A vssd1 vssd1 vccd1 vccd1 _20980_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19639_ _19639_/A vssd1 vssd1 vccd1 vccd1 _19639_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22650_ _22698_/A vssd1 vssd1 vccd1 vccd1 _22650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21601_ _21649_/A vssd1 vssd1 vccd1 vccd1 _21601_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22581_ _22597_/A vssd1 vssd1 vccd1 vccd1 _22581_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24320_ _27544_/Q _24328_/B vssd1 vssd1 vccd1 vccd1 _24321_/A sky130_fd_sc_hd__and2_1
X_21532_ _21564_/A vssd1 vssd1 vccd1 vccd1 _21532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24251_ _24251_/A vssd1 vssd1 vccd1 vccd1 _27397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21463_ _21463_/A vssd1 vssd1 vccd1 vccd1 _21463_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23202_ _17450_/X _27138_/Q _23204_/S vssd1 vssd1 vccd1 vccd1 _23203_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20414_ _20408_/X _20409_/X _20410_/X _20411_/X _20412_/X _20413_/X vssd1 vssd1 vccd1
+ vccd1 _20415_/A sky130_fd_sc_hd__mux4_1
X_24182_ _27467_/Q _24184_/B vssd1 vssd1 vccd1 vccd1 _24183_/A sky130_fd_sc_hd__and2_1
XFILLER_105_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21394_ _21463_/A vssd1 vssd1 vccd1 vccd1 _21394_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23133_ _23133_/A vssd1 vssd1 vccd1 vccd1 _27107_/D sky130_fd_sc_hd__clkbuf_1
X_20345_ _20345_/A vssd1 vssd1 vccd1 vccd1 _20345_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23064_ _27077_/Q _17712_/X _23070_/S vssd1 vssd1 vccd1 vccd1 _23065_/A sky130_fd_sc_hd__mux2_1
X_27941_ _27941_/A _15941_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
X_20276_ _20267_/X _20269_/X _20271_/X _20273_/X _20274_/X _20275_/X vssd1 vssd1 vccd1
+ vccd1 _20277_/A sky130_fd_sc_hd__mux4_1
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22015_ _22015_/A vssd1 vssd1 vccd1 vccd1 _22083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26823_ _22190_/X _26823_/D vssd1 vssd1 vccd1 vccd1 _26823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26754_ _21948_/X _26754_/D vssd1 vssd1 vccd1 vccd1 _26754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23966_ _23943_/X _23964_/X _23965_/X _23958_/X vssd1 vssd1 vccd1 vccd1 _27292_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25705_ _25721_/A vssd1 vssd1 vccd1 vccd1 _25705_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22917_ _22907_/X _22908_/X _22909_/X _22910_/X _22911_/X _22912_/X vssd1 vssd1 vccd1
+ vccd1 _22918_/A sky130_fd_sc_hd__mux4_1
XFILLER_99_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23897_ _23991_/A vssd1 vssd1 vccd1 vccd1 _23897_/X sky130_fd_sc_hd__clkbuf_2
X_26685_ _21712_/X _26685_/D vssd1 vssd1 vccd1 vccd1 _26685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13650_ _13921_/A _13661_/B vssd1 vssd1 vccd1 vccd1 _13650_/Y sky130_fd_sc_hd__nor2_1
X_22848_ _22848_/A vssd1 vssd1 vccd1 vccd1 _22848_/X sky130_fd_sc_hd__clkbuf_1
X_25636_ _25636_/A vssd1 vssd1 vccd1 vccd1 _25636_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13581_ _27335_/Q _13022_/X _13030_/X _27303_/Q _13237_/X vssd1 vssd1 vccd1 vccd1
+ _14531_/A sky130_fd_sc_hd__a221oi_4
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25567_ _25560_/X _25291_/B _25565_/X _25566_/X vssd1 vssd1 vccd1 vccd1 _25567_/X
+ sky130_fd_sc_hd__a211o_1
X_22779_ _22767_/X _22768_/X _22769_/X _22770_/X _22771_/X _22772_/X vssd1 vssd1 vccd1
+ vccd1 _22780_/A sky130_fd_sc_hd__mux4_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15320_ _26304_/Q _13401_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__mux2_1
X_27306_ _27379_/CLK _27306_/D vssd1 vssd1 vccd1 vccd1 _27306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24518_ _24518_/A vssd1 vssd1 vccd1 vccd1 _27528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25498_ _24759_/A _25474_/X _25491_/Y _25496_/X _25497_/X vssd1 vssd1 vccd1 vccd1
+ _27763_/D sky130_fd_sc_hd__a221oi_1
XFILLER_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15251_ _15251_/A vssd1 vssd1 vccd1 vccd1 _26335_/D sky130_fd_sc_hd__clkbuf_1
X_27237_ _27264_/CLK _27237_/D vssd1 vssd1 vccd1 vccd1 _27237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24449_ _24449_/A vssd1 vssd1 vccd1 vccd1 _27501_/D sky130_fd_sc_hd__clkbuf_1
X_14202_ _14215_/A vssd1 vssd1 vccd1 vccd1 _14213_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15182_ _26365_/Q _13411_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27168_ _27225_/CLK _27168_/D vssd1 vssd1 vccd1 vccd1 _27168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14133_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14133_/X sky130_fd_sc_hd__clkbuf_2
X_26119_ _19725_/X _26119_/D vssd1 vssd1 vccd1 vccd1 _26119_/Q sky130_fd_sc_hd__dfxtp_1
X_19990_ _19990_/A vssd1 vssd1 vccd1 vccd1 _19990_/X sky130_fd_sc_hd__clkbuf_1
X_27099_ _27410_/CLK _27099_/D vssd1 vssd1 vccd1 vccd1 _27099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ _14147_/B vssd1 vssd1 vccd1 vccd1 _14064_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18941_ _19387_/A vssd1 vssd1 vccd1 vccd1 _18941_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ _27367_/Q _27368_/Q vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__and2b_1
XFILLER_106_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18872_ _18969_/A _18872_/B vssd1 vssd1 vccd1 vccd1 _18872_/X sky130_fd_sc_hd__or2_1
XFILLER_79_465 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17823_ _18403_/A vssd1 vssd1 vccd1 vccd1 _17959_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17754_ _25936_/Q _17753_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17755_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14966_ _15703_/A _14966_/B vssd1 vssd1 vccd1 vccd1 _14966_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16705_ _16744_/A _16372_/A _16704_/X vssd1 vssd1 vccd1 vccd1 _16705_/X sky130_fd_sc_hd__o21a_1
X_13917_ _13917_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _13917_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17685_ _17685_/A vssd1 vssd1 vccd1 vccd1 _25914_/D sky130_fd_sc_hd__clkbuf_1
X_14897_ _14897_/A vssd1 vssd1 vccd1 vccd1 _26485_/D sky130_fd_sc_hd__clkbuf_1
X_19424_ _19422_/X _19423_/X _19468_/S vssd1 vssd1 vccd1 vccd1 _19424_/X sky130_fd_sc_hd__mux2_2
X_16636_ _16584_/Y _16636_/B vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__and2b_1
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13848_ _26842_/Q _13844_/X _13770_/B _13847_/Y vssd1 vssd1 vccd1 vccd1 _26842_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_16_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28009__475 vssd1 vssd1 vccd1 vccd1 _28009__475/HI _28009_/A sky130_fd_sc_hd__conb_1
X_19355_ _19351_/X _19353_/X _19354_/X vssd1 vssd1 vccd1 vccd1 _19355_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16567_ _16798_/A _16567_/B vssd1 vssd1 vccd1 vccd1 _16572_/B sky130_fd_sc_hd__xor2_1
X_13779_ _13779_/A vssd1 vssd1 vccd1 vccd1 _13833_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18306_ _26412_/Q _26380_/Q _26348_/Q _26316_/Q _18305_/X _18214_/X vssd1 vssd1 vccd1
+ vccd1 _18306_/X sky130_fd_sc_hd__mux4_1
X_15518_ _15518_/A vssd1 vssd1 vccd1 vccd1 _26217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19286_ _26412_/Q _26380_/Q _26348_/Q _26316_/Q _19170_/X _19240_/X vssd1 vssd1 vccd1
+ vccd1 _19286_/X sky130_fd_sc_hd__mux4_1
X_16498_ _16499_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16500_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18237_ _18234_/X _18235_/X _18331_/S vssd1 vssd1 vccd1 vccd1 _18237_/X sky130_fd_sc_hd__mux2_1
X_15449_ _26247_/Q _13379_/X _15451_/S vssd1 vssd1 vccd1 vccd1 _15450_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1069 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18168_ _18285_/A vssd1 vssd1 vccd1 vccd1 _18168_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17119_ _17094_/X _17119_/B vssd1 vssd1 vccd1 vccd1 _17119_/X sky130_fd_sc_hd__and2b_1
X_18099_ _18401_/A vssd1 vssd1 vccd1 vccd1 _18099_/X sky130_fd_sc_hd__buf_2
XFILLER_132_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20130_ _20162_/A vssd1 vssd1 vccd1 vccd1 _20130_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20061_ _20077_/A vssd1 vssd1 vccd1 vccd1 _20061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater220 _27401_/CLK vssd1 vssd1 vccd1 vccd1 _27398_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater231 _26062_/CLK vssd1 vssd1 vccd1 vccd1 _26069_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater242 _27606_/CLK vssd1 vssd1 vccd1 vccd1 _27752_/CLK sky130_fd_sc_hd__clkbuf_1
X_23820_ _23818_/X _23819_/X _23844_/S vssd1 vssd1 vccd1 vccd1 _23820_/X sky130_fd_sc_hd__mux2_1
Xrepeater253 _27621_/CLK vssd1 vssd1 vccd1 vccd1 _27700_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater264 _27185_/CLK vssd1 vssd1 vccd1 vccd1 _27180_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater275 _27539_/CLK vssd1 vssd1 vccd1 vccd1 _27534_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23751_ _27787_/Q vssd1 vssd1 vccd1 vccd1 _24045_/S sky130_fd_sc_hd__buf_2
Xrepeater286 _27372_/CLK vssd1 vssd1 vccd1 vccd1 _27480_/CLK sky130_fd_sc_hd__clkbuf_1
XANTENNA_309 _18079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20963_ _20953_/X _20954_/X _20955_/X _20956_/X _20958_/X _20960_/X vssd1 vssd1 vccd1
+ vccd1 _20964_/A sky130_fd_sc_hd__mux4_1
Xrepeater297 _27264_/CLK vssd1 vssd1 vccd1 vccd1 _27263_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22702_ _22771_/A vssd1 vssd1 vccd1 vccd1 _22702_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23682_ _23682_/A vssd1 vssd1 vccd1 vccd1 _27246_/D sky130_fd_sc_hd__clkbuf_1
X_26470_ _20962_/X _26470_/D vssd1 vssd1 vccd1 vccd1 _26470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20894_ _20942_/A vssd1 vssd1 vccd1 vccd1 _20894_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22633_ _22891_/A vssd1 vssd1 vccd1 vccd1 _22699_/A sky130_fd_sc_hd__buf_2
X_25421_ _25421_/A vssd1 vssd1 vccd1 vccd1 _27748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25352_ _27719_/Q _25139_/A _25351_/Y _13423_/X vssd1 vssd1 vccd1 vccd1 _27719_/D
+ sky130_fd_sc_hd__o211a_1
X_22564_ _22612_/A vssd1 vssd1 vccd1 vccd1 _22564_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21515_ _21563_/A vssd1 vssd1 vccd1 vccd1 _21515_/X sky130_fd_sc_hd__clkbuf_1
X_24303_ _16296_/X _16297_/Y _16298_/X _24217_/A vssd1 vssd1 vccd1 vccd1 _27433_/D
+ sky130_fd_sc_hd__a31oi_4
XFILLER_22_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25283_ _25306_/A _25283_/B vssd1 vssd1 vccd1 vccd1 _25283_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22495_ _22487_/X _22488_/X _22489_/X _22490_/X _22491_/X _22492_/X vssd1 vssd1 vccd1
+ vccd1 _22496_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27022_ _22882_/X _27022_/D vssd1 vssd1 vccd1 vccd1 _27022_/Q sky130_fd_sc_hd__dfxtp_1
X_24234_ _24234_/A vssd1 vssd1 vccd1 vccd1 _27388_/D sky130_fd_sc_hd__clkbuf_1
X_21446_ _21478_/A vssd1 vssd1 vccd1 vccd1 _21446_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24165_ _27459_/Q _24173_/B vssd1 vssd1 vccd1 vccd1 _24166_/A sky130_fd_sc_hd__and2_1
X_21377_ _21377_/A vssd1 vssd1 vccd1 vccd1 _21377_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23116_ _23116_/A vssd1 vssd1 vccd1 vccd1 _27099_/D sky130_fd_sc_hd__clkbuf_1
X_20328_ _20318_/X _20319_/X _20320_/X _20321_/X _20322_/X _20323_/X vssd1 vssd1 vccd1
+ vccd1 _20329_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24096_ _24096_/A vssd1 vssd1 vccd1 vccd1 _27323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27924_ _27924_/A _15963_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
X_23047_ _23047_/A vssd1 vssd1 vccd1 vccd1 _27069_/D sky130_fd_sc_hd__clkbuf_1
X_20259_ _20259_/A vssd1 vssd1 vccd1 vccd1 _20259_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27855_ _27855_/CLK _27855_/D vssd1 vssd1 vccd1 vccd1 _27855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26806_ _22134_/X _26806_/D vssd1 vssd1 vccd1 vccd1 _26806_/Q sky130_fd_sc_hd__dfxtp_1
X_14820_ _26519_/Q _13328_/X _14824_/S vssd1 vssd1 vccd1 vccd1 _14821_/A sky130_fd_sc_hd__mux2_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27786_ _27786_/CLK _27786_/D vssd1 vssd1 vccd1 vccd1 _27786_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24998_ _24994_/X _24995_/X _25031_/S vssd1 vssd1 vccd1 vccd1 _24998_/X sky130_fd_sc_hd__mux2_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26737_ _21890_/X _26737_/D vssd1 vssd1 vccd1 vccd1 _26737_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14750_/X _26541_/Q _14757_/S vssd1 vssd1 vccd1 vccd1 _14752_/A sky130_fd_sc_hd__mux2_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23949_ _23945_/X _23947_/X _23985_/S vssd1 vssd1 vccd1 vccd1 _23949_/X sky130_fd_sc_hd__mux2_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _26897_/Q _13697_/X _13692_/X _13701_/Y vssd1 vssd1 vccd1 vccd1 _26897_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17470_ _17469_/X _25825_/Q _17470_/S vssd1 vssd1 vccd1 vccd1 _17471_/A sky130_fd_sc_hd__mux2_1
X_26668_ _21644_/X _26668_/D vssd1 vssd1 vccd1 vccd1 _26668_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _15756_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14682_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16421_ _14775_/A _16314_/X _16098_/A _25955_/Q _16420_/Y vssd1 vssd1 vccd1 vccd1
+ _16772_/B sky130_fd_sc_hd__a221o_1
X_13633_ _26921_/Q _13626_/X _13629_/X _13632_/Y vssd1 vssd1 vccd1 vccd1 _26921_/D
+ sky130_fd_sc_hd__a31o_1
X_25619_ _23638_/A _27979_/A _25623_/S vssd1 vssd1 vccd1 vccd1 _25620_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26599_ _21406_/X _26599_/D vssd1 vssd1 vccd1 vccd1 _26599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19140_ _18895_/X _19134_/X _19136_/X _19138_/X _19139_/X vssd1 vssd1 vccd1 vccd1
+ _19153_/B sky130_fd_sc_hd__a221o_1
X_16352_ _16332_/X _16858_/B _16857_/A vssd1 vssd1 vccd1 vccd1 _16674_/A sky130_fd_sc_hd__a21oi_1
XFILLER_198_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13564_ _14518_/A vssd1 vssd1 vccd1 vccd1 _13930_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_197_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ _15303_/A vssd1 vssd1 vccd1 vccd1 _26312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19071_ _26147_/Q _26083_/Q _27011_/Q _26979_/Q _19049_/X _19070_/X vssd1 vssd1 vccd1
+ vccd1 _19072_/B sky130_fd_sc_hd__mux4_1
X_13495_ _26957_/Q _13487_/X _13482_/X _13494_/Y vssd1 vssd1 vccd1 vccd1 _26957_/D
+ sky130_fd_sc_hd__a31o_1
X_16283_ _27396_/Q _16298_/B vssd1 vssd1 vccd1 vccd1 _16283_/Y sky130_fd_sc_hd__nand2_1
XFILLER_201_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18022_ _18020_/X _18021_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _18022_/X sky130_fd_sc_hd__o21a_1
X_15234_ _14772_/X _26342_/Q _15234_/S vssd1 vssd1 vccd1 vccd1 _15235_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1080 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15165_ _26373_/Q _13385_/X _15173_/S vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _26759_/Q _14104_/X _14107_/X _14115_/Y vssd1 vssd1 vccd1 vccd1 _26759_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ _15096_/A vssd1 vssd1 vccd1 vccd1 _26404_/D sky130_fd_sc_hd__clkbuf_1
X_19973_ _19989_/A vssd1 vssd1 vccd1 vccd1 _19973_/X sky130_fd_sc_hd__clkbuf_1
X_18924_ _26525_/Q _26493_/Q _26461_/Q _27037_/Q _18922_/X _18923_/X vssd1 vssd1 vccd1
+ vccd1 _18924_/X sky130_fd_sc_hd__mux4_1
X_14047_ _14403_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18855_ _18846_/X _18849_/X _18853_/X _18854_/X _24407_/A vssd1 vssd1 vccd1 vccd1
+ _18868_/B sky130_fd_sc_hd__a221o_1
XFILLER_68_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17806_ _26810_/Q _26778_/Q _26746_/Q _26714_/Q _17801_/X _17805_/X vssd1 vssd1 vccd1
+ vccd1 _17806_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18786_ _18775_/X _18783_/X _18785_/X vssd1 vssd1 vccd1 vccd1 _18786_/X sky130_fd_sc_hd__o21a_1
X_15998_ _27481_/Q _27372_/Q vssd1 vssd1 vccd1 vccd1 _16001_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17737_ _27427_/Q vssd1 vssd1 vccd1 vccd1 _17737_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14949_ _14801_/X _26461_/Q _14951_/S vssd1 vssd1 vccd1 vccd1 _14950_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17668_ _17668_/A vssd1 vssd1 vccd1 vccd1 _25904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19407_ _19407_/A vssd1 vssd1 vccd1 vccd1 _19407_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16619_ _16619_/A vssd1 vssd1 vccd1 vccd1 _16619_/X sky130_fd_sc_hd__clkbuf_2
X_17599_ _17523_/X _25874_/Q _17599_/S vssd1 vssd1 vccd1 vccd1 _17600_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19338_ _19338_/A vssd1 vssd1 vccd1 vccd1 _19338_/X sky130_fd_sc_hd__buf_2
XFILLER_148_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19269_ _19269_/A vssd1 vssd1 vccd1 vccd1 _26059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_191_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21300_ _21300_/A vssd1 vssd1 vccd1 vccd1 _21300_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22280_ _22347_/A vssd1 vssd1 vccd1 vccd1 _22280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21231_ _21301_/A vssd1 vssd1 vccd1 vccd1 _21231_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21162_ _21162_/A vssd1 vssd1 vccd1 vccd1 _21162_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20113_ _20113_/A vssd1 vssd1 vccd1 vccd1 _20113_/X sky130_fd_sc_hd__clkbuf_1
X_25970_ _25974_/CLK _25970_/D vssd1 vssd1 vccd1 vccd1 _25970_/Q sky130_fd_sc_hd__dfxtp_1
X_21093_ _21125_/A vssd1 vssd1 vccd1 vccd1 _21093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20044_ _20076_/A vssd1 vssd1 vccd1 vccd1 _20044_/X sky130_fd_sc_hd__clkbuf_1
X_24921_ _27660_/Q _24909_/X _24920_/Y _24914_/X vssd1 vssd1 vccd1 vccd1 _27660_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27640_ _27690_/CLK _27640_/D vssd1 vssd1 vccd1 vccd1 _27640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24852_ _24848_/A _24851_/C _27760_/Q vssd1 vssd1 vccd1 vccd1 _24853_/B sky130_fd_sc_hd__a21oi_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23803_ _27831_/Q _27135_/Q _25880_/Q _25848_/Q _23777_/X _23802_/X vssd1 vssd1 vccd1
+ vccd1 _23803_/X sky130_fd_sc_hd__mux4_1
X_27571_ _27575_/CLK _27571_/D vssd1 vssd1 vccd1 vccd1 _27571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _21981_/X _21982_/X _21983_/X _21984_/X _21985_/X _21986_/X vssd1 vssd1 vccd1
+ vccd1 _21996_/A sky130_fd_sc_hd__mux4_1
XFILLER_22_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24783_ _27627_/Q _24771_/X _24782_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _27627_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_1136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_106 _19519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _22540_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_128 _20942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26522_ _21138_/X _26522_/D vssd1 vssd1 vccd1 vccd1 _26522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _15773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20946_ _20946_/A vssd1 vssd1 vccd1 vccd1 _20946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23734_ _27373_/Q _24050_/B vssd1 vssd1 vccd1 vccd1 _23735_/A sky130_fd_sc_hd__and2_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26453_ _20902_/X _26453_/D vssd1 vssd1 vccd1 vccd1 _26453_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20877_ _20864_/X _20865_/X _20866_/X _20867_/X _20870_/X _20874_/X vssd1 vssd1 vccd1
+ vccd1 _20878_/A sky130_fd_sc_hd__mux4_1
X_23665_ _23665_/A vssd1 vssd1 vccd1 vccd1 _27238_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25404_ _25415_/A vssd1 vssd1 vccd1 vccd1 _25413_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22616_ _22616_/A vssd1 vssd1 vccd1 vccd1 _22961_/A sky130_fd_sc_hd__buf_2
X_23596_ _23596_/A _23596_/B vssd1 vssd1 vccd1 vccd1 _23597_/A sky130_fd_sc_hd__and2_1
X_26384_ _20651_/X _26384_/D vssd1 vssd1 vccd1 vccd1 _26384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22547_ _22893_/A vssd1 vssd1 vccd1 vccd1 _22612_/A sky130_fd_sc_hd__buf_2
X_25335_ _25339_/B _25335_/B vssd1 vssd1 vccd1 vccd1 _25336_/B sky130_fd_sc_hd__nand2_1
XFILLER_167_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13280_ _27019_/Q _13139_/X _13280_/S vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__mux2_1
X_22478_ _22478_/A vssd1 vssd1 vccd1 vccd1 _22478_/X sky130_fd_sc_hd__clkbuf_1
X_25266_ _25266_/A _25266_/B _25242_/B _25265_/Y vssd1 vssd1 vccd1 vccd1 _25272_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_136_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27005_ _22828_/X _27005_/D vssd1 vssd1 vccd1 vccd1 _27005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21429_ _21477_/A vssd1 vssd1 vccd1 vccd1 _21429_/X sky130_fd_sc_hd__clkbuf_1
X_24217_ _24217_/A vssd1 vssd1 vccd1 vccd1 _24222_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25197_ _25197_/A _25197_/B vssd1 vssd1 vccd1 vccd1 _25198_/B sky130_fd_sc_hd__nand2_1
XFILLER_151_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24148_ _24148_/A vssd1 vssd1 vccd1 vccd1 _27346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16970_ _24435_/A vssd1 vssd1 vccd1 vccd1 _24636_/A sky130_fd_sc_hd__clkbuf_1
X_24079_ _24079_/A vssd1 vssd1 vccd1 vccd1 _27315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15921_ _15924_/A vssd1 vssd1 vccd1 vccd1 _15921_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18640_ _18640_/A vssd1 vssd1 vccd1 vccd1 _25986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27838_ _27840_/CLK _27838_/D vssd1 vssd1 vccd1 vccd1 _27838_/Q sky130_fd_sc_hd__dfxtp_1
X_15852_ _15852_/A vssd1 vssd1 vccd1 vccd1 _26075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14803_/A vssd1 vssd1 vccd1 vccd1 _26525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _18571_/A _18474_/X vssd1 vssd1 vccd1 vccd1 _18571_/X sky130_fd_sc_hd__or2b_1
XFILLER_18_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27769_ _27774_/CLK _27769_/D vssd1 vssd1 vccd1 vccd1 _27769_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15783_ _15783_/A _15783_/B vssd1 vssd1 vccd1 vccd1 _15840_/A sky130_fd_sc_hd__or2_2
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _12995_/A vssd1 vssd1 vccd1 vccd1 _27801_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _17522_/A vssd1 vssd1 vccd1 vccd1 _25841_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14734_ _14734_/A vssd1 vssd1 vccd1 vccd1 _14734_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_189_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _27417_/Q vssd1 vssd1 vccd1 vccd1 _17453_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14665_ _26571_/Q _14658_/X _14653_/X _14664_/Y vssd1 vssd1 vccd1 vccd1 _26571_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16404_ _14500_/A _16563_/B _16067_/X _16401_/Y _16403_/Y vssd1 vssd1 vccd1 vccd1
+ _16774_/B sky130_fd_sc_hd__o221a_1
XFILLER_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ _13656_/A vssd1 vssd1 vccd1 vccd1 _13616_/X sky130_fd_sc_hd__clkbuf_2
X_17384_ _17116_/A _17379_/X _17381_/X _17383_/X vssd1 vssd1 vccd1 vccd1 _17384_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_186_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14596_ _26596_/Q _14589_/X _14592_/X _14595_/Y vssd1 vssd1 vccd1 vccd1 _26596_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19123_ _19123_/A _19123_/B vssd1 vssd1 vccd1 vccd1 _19123_/X sky130_fd_sc_hd__or2_1
XFILLER_71_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16335_ _16756_/B vssd1 vssd1 vccd1 vccd1 _16753_/B sky130_fd_sc_hd__clkbuf_1
X_13547_ _13921_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13547_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19054_ _19343_/A vssd1 vssd1 vccd1 vccd1 _19054_/X sky130_fd_sc_hd__buf_2
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16266_ _16266_/A _27535_/Q vssd1 vssd1 vccd1 vccd1 _16266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13478_ _27357_/Q _13021_/A _13102_/X _27325_/Q _13109_/X vssd1 vssd1 vccd1 vccd1
+ _14452_/A sky130_fd_sc_hd__a221oi_4
X_18005_ _18481_/A vssd1 vssd1 vccd1 vccd1 _18005_/X sky130_fd_sc_hd__clkbuf_2
X_15217_ _14747_/X _26350_/Q _15223_/S vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16197_ _16197_/A _16215_/B _16197_/C vssd1 vssd1 vccd1 vccd1 _16197_/X sky130_fd_sc_hd__and3_1
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15148_ _15148_/A vssd1 vssd1 vccd1 vccd1 _26381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15079_ _14756_/X _26411_/Q _15079_/S vssd1 vssd1 vccd1 vccd1 _15080_/A sky130_fd_sc_hd__mux2_1
X_19956_ _19988_/A vssd1 vssd1 vccd1 vccd1 _19956_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18907_ _18922_/A vssd1 vssd1 vccd1 vccd1 _19441_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19887_ _19887_/A vssd1 vssd1 vccd1 vccd1 _19887_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18838_ _27602_/Q vssd1 vssd1 vccd1 vccd1 _19469_/A sky130_fd_sc_hd__inv_2
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18769_ _19460_/A vssd1 vssd1 vccd1 vccd1 _19486_/A sky130_fd_sc_hd__buf_2
X_20800_ _20800_/A vssd1 vssd1 vccd1 vccd1 _22546_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21780_ _21828_/A vssd1 vssd1 vccd1 vccd1 _21780_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20731_ _20731_/A vssd1 vssd1 vccd1 vccd1 _20731_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23450_ input11/X _23442_/X _23449_/X _23447_/X vssd1 vssd1 vccd1 vccd1 _27173_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20662_ _20652_/X _20653_/X _20654_/X _20655_/X _20656_/X _20657_/X vssd1 vssd1 vccd1
+ vccd1 _20663_/A sky130_fd_sc_hd__mux4_1
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22401_ _22433_/A vssd1 vssd1 vccd1 vccd1 _22401_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23381_ _27756_/Q _23376_/Y _27240_/Q _24752_/A _23380_/X vssd1 vssd1 vccd1 vccd1
+ _23393_/A sky130_fd_sc_hd__a221o_1
X_20593_ _20593_/A vssd1 vssd1 vccd1 vccd1 _20593_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22332_ _22348_/A vssd1 vssd1 vccd1 vccd1 _22332_/X sky130_fd_sc_hd__clkbuf_1
X_25120_ _27521_/Q _27489_/Q vssd1 vssd1 vccd1 vccd1 _25129_/A sky130_fd_sc_hd__or2_1
XFILLER_191_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25051_ _27835_/Q _27139_/Q _25884_/Q _25852_/Q _25018_/X _25035_/X vssd1 vssd1 vccd1
+ vccd1 _25051_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22263_ _22263_/A vssd1 vssd1 vccd1 vccd1 _22263_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24002_ _24002_/A vssd1 vssd1 vccd1 vccd1 _24002_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21214_ _21214_/A vssd1 vssd1 vccd1 vccd1 _21214_/X sky130_fd_sc_hd__clkbuf_1
X_22194_ _22261_/A vssd1 vssd1 vccd1 vccd1 _22194_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21145_ _21145_/A vssd1 vssd1 vccd1 vccd1 _21212_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_487 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21076_ _21076_/A vssd1 vssd1 vccd1 vccd1 _21076_/X sky130_fd_sc_hd__clkbuf_1
X_25953_ _25953_/CLK _25953_/D vssd1 vssd1 vccd1 vccd1 _25953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24904_ _24913_/A _24904_/B vssd1 vssd1 vccd1 vccd1 _24904_/Y sky130_fd_sc_hd__nand2_1
X_20027_ _20027_/A vssd1 vssd1 vccd1 vccd1 _20027_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25884_ _25884_/CLK _25884_/D vssd1 vssd1 vccd1 vccd1 _25884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27623_ _27623_/CLK _27623_/D vssd1 vssd1 vccd1 vccd1 _27623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24835_ _24835_/A _24835_/B _27755_/Q vssd1 vssd1 vccd1 vccd1 _24844_/B sky130_fd_sc_hd__and3_1
XFILLER_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27554_ _27558_/CLK _27554_/D vssd1 vssd1 vccd1 vccd1 _27554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24766_ _27620_/Q _24758_/X _24765_/Y _24760_/X vssd1 vssd1 vccd1 vccd1 _27620_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _21978_/A vssd1 vssd1 vccd1 vccd1 _21978_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26505_ _21084_/X _26505_/D vssd1 vssd1 vccd1 vccd1 _26505_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23717_ _23717_/A vssd1 vssd1 vccd1 vccd1 _27262_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20929_ _20921_/X _20922_/X _20923_/X _20924_/X _20925_/X _20926_/X vssd1 vssd1 vccd1
+ vccd1 _20930_/A sky130_fd_sc_hd__mux4_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27485_ _27600_/CLK _27485_/D vssd1 vssd1 vccd1 vccd1 _27485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24697_ _24394_/A _24687_/X _24696_/X _24690_/X vssd1 vssd1 vccd1 vccd1 _27596_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _15723_/A _14465_/B vssd1 vssd1 vccd1 vccd1 _14450_/Y sky130_fd_sc_hd__nor2_1
X_26436_ _20841_/X _26436_/D vssd1 vssd1 vccd1 vccd1 _26436_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23648_ _23643_/X _24987_/S _23638_/X _25623_/S vssd1 vssd1 vccd1 vccd1 _23649_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13401_ _14791_/A vssd1 vssd1 vccd1 vccd1 _13401_/X sky130_fd_sc_hd__clkbuf_4
X_14381_ _14381_/A _14390_/B vssd1 vssd1 vccd1 vccd1 _14381_/Y sky130_fd_sc_hd__nor2_1
X_26367_ _20593_/X _26367_/D vssd1 vssd1 vccd1 vccd1 _26367_/Q sky130_fd_sc_hd__dfxtp_1
X_23579_ _23598_/A vssd1 vssd1 vccd1 vccd1 _23596_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16120_ _16252_/B _16252_/C vssd1 vssd1 vccd1 vccd1 _16277_/B sky130_fd_sc_hd__nand2_2
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25318_ _25319_/B _25319_/C _25328_/A vssd1 vssd1 vccd1 vccd1 _25320_/A sky130_fd_sc_hd__a21oi_1
X_13332_ _26998_/Q _13331_/X _13335_/S vssd1 vssd1 vccd1 vccd1 _13333_/A sky130_fd_sc_hd__mux2_1
X_26298_ _20349_/X _26298_/D vssd1 vssd1 vccd1 vccd1 _26298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ _16066_/A _16066_/B _16066_/C vssd1 vssd1 vccd1 vccd1 _16353_/A sky130_fd_sc_hd__nand3_2
XFILLER_143_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25249_ _25249_/A _25267_/A vssd1 vssd1 vccd1 vccd1 _25265_/A sky130_fd_sc_hd__nand2_1
X_13263_ _27027_/Q _13094_/X _13269_/S vssd1 vssd1 vccd1 vccd1 _13264_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15002_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13194_ _13194_/A vssd1 vssd1 vccd1 vccd1 _13194_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19810_ _19796_/X _19797_/X _19798_/X _19799_/X _19800_/X _19801_/X vssd1 vssd1 vccd1
+ vccd1 _19811_/A sky130_fd_sc_hd__mux4_1
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19741_ _19741_/A vssd1 vssd1 vccd1 vccd1 _19741_/X sky130_fd_sc_hd__clkbuf_1
X_16953_ _27583_/Q vssd1 vssd1 vccd1 vccd1 _24635_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15904_ _15906_/A vssd1 vssd1 vccd1 vccd1 _15904_/Y sky130_fd_sc_hd__inv_2
X_19672_ _19659_/X _19661_/X _19663_/X _19665_/X _19666_/X _19667_/X vssd1 vssd1 vccd1
+ vccd1 _19673_/A sky130_fd_sc_hd__mux4_1
X_16884_ _16077_/X _16802_/A _16616_/A _16650_/A vssd1 vssd1 vccd1 vccd1 _16884_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18623_ _18623_/A vssd1 vssd1 vccd1 vccd1 _25978_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _15835_/A vssd1 vssd1 vccd1 vccd1 _26083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18554_ _18009_/X _18551_/X _18553_/X _18014_/X vssd1 vssd1 vccd1 vccd1 _18554_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15766_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12978_ _13000_/A vssd1 vssd1 vccd1 vccd1 _12987_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17505_ _17505_/A vssd1 vssd1 vccd1 vccd1 _17518_/S sky130_fd_sc_hd__buf_2
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _14717_/A vssd1 vssd1 vccd1 vccd1 _26552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18485_ _26548_/Q _26516_/Q _26484_/Q _27060_/Q _18392_/X _18418_/X vssd1 vssd1 vccd1
+ vccd1 _18485_/X sky130_fd_sc_hd__mux4_1
X_15697_ _15781_/B vssd1 vssd1 vccd1 vccd1 _15697_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17436_ _17436_/A vssd1 vssd1 vccd1 vccd1 _25814_/D sky130_fd_sc_hd__clkbuf_1
X_14648_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14659_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_17 _25992_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _27296_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_39 _17898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _27224_/Q _17366_/X _17367_/S vssd1 vssd1 vccd1 vccd1 _17368_/A sky130_fd_sc_hd__mux2_1
X_14579_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14579_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19106_ _19097_/X _19099_/X _19104_/X _19035_/X _19105_/X vssd1 vssd1 vccd1 vccd1
+ _19107_/C sky130_fd_sc_hd__a221o_1
XFILLER_192_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16318_ _16593_/B _16595_/B _16639_/A vssd1 vssd1 vccd1 vccd1 _16319_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17298_ _17298_/A vssd1 vssd1 vccd1 vccd1 _27939_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19037_ _19107_/A _19037_/B _19037_/C vssd1 vssd1 vccd1 vccd1 _19038_/A sky130_fd_sc_hd__and3_1
X_16249_ _16249_/A _16249_/B _16252_/C vssd1 vssd1 vccd1 vccd1 _16249_/X sky130_fd_sc_hd__and3_1
XFILLER_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19939_ _19939_/A vssd1 vssd1 vccd1 vccd1 _19939_/X sky130_fd_sc_hd__clkbuf_1
X_22950_ _22950_/A vssd1 vssd1 vccd1 vccd1 _22950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21901_ _21895_/X _21896_/X _21897_/X _21898_/X _21899_/X _21900_/X vssd1 vssd1 vccd1
+ vccd1 _21902_/A sky130_fd_sc_hd__mux4_1
X_22881_ _22869_/X _22870_/X _22871_/X _22872_/X _22874_/X _22876_/X vssd1 vssd1 vccd1
+ vccd1 _22882_/A sky130_fd_sc_hd__mux4_1
XFILLER_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24620_ _27669_/Q _24620_/B vssd1 vssd1 vccd1 vccd1 _24621_/A sky130_fd_sc_hd__and2_1
X_21832_ _21900_/A vssd1 vssd1 vccd1 vccd1 _21832_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21763_ _22021_/A vssd1 vssd1 vccd1 vccd1 _21828_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24551_ _27609_/Q _18352_/S _24551_/S vssd1 vssd1 vccd1 vccd1 _24552_/B sky130_fd_sc_hd__mux2_1
XFILLER_168_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20714_ _20703_/X _20705_/X _20707_/X _20709_/X _20710_/X _20711_/X vssd1 vssd1 vccd1
+ vccd1 _20715_/A sky130_fd_sc_hd__mux4_2
X_23502_ input8/X input7/X vssd1 vssd1 vccd1 vccd1 _23650_/B sky130_fd_sc_hd__and2_4
XFILLER_93_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27270_ _27335_/CLK _27270_/D vssd1 vssd1 vccd1 vccd1 _27270_/Q sky130_fd_sc_hd__dfxtp_2
X_21694_ _21726_/A vssd1 vssd1 vccd1 vccd1 _21694_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24482_ _24482_/A vssd1 vssd1 vccd1 vccd1 _27516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26221_ _20087_/X _26221_/D vssd1 vssd1 vccd1 vccd1 _26221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20645_ _20645_/A vssd1 vssd1 vccd1 vccd1 _20645_/X sky130_fd_sc_hd__clkbuf_1
X_23433_ _27167_/Q _23443_/B vssd1 vssd1 vccd1 vccd1 _23433_/X sky130_fd_sc_hd__or2_1
XFILLER_184_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23364_ _27771_/Q vssd1 vssd1 vccd1 vccd1 _24906_/A sky130_fd_sc_hd__buf_4
X_26152_ _19845_/X _26152_/D vssd1 vssd1 vccd1 vccd1 _26152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20576_ _20566_/X _20567_/X _20568_/X _20569_/X _20570_/X _20571_/X vssd1 vssd1 vccd1
+ vccd1 _20577_/A sky130_fd_sc_hd__mux4_1
XFILLER_137_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25103_ _25101_/X _25102_/X _25103_/S vssd1 vssd1 vccd1 vccd1 _25103_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22315_ _22347_/A vssd1 vssd1 vccd1 vccd1 _22315_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23295_ input47/X vssd1 vssd1 vccd1 vccd1 _23295_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26083_ _19602_/X _26083_/D vssd1 vssd1 vccd1 vccd1 _26083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22246_ _22262_/A vssd1 vssd1 vccd1 vccd1 _22246_/X sky130_fd_sc_hd__clkbuf_1
X_25034_ _25034_/A vssd1 vssd1 vccd1 vccd1 _27678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22177_ _22613_/A vssd1 vssd1 vccd1 vccd1 _22523_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21128_ _21128_/A vssd1 vssd1 vccd1 vccd1 _21128_/X sky130_fd_sc_hd__clkbuf_1
X_26985_ _22758_/X _26985_/D vssd1 vssd1 vccd1 vccd1 _26985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25936_ _27124_/CLK _25936_/D vssd1 vssd1 vccd1 vccd1 _25936_/Q sky130_fd_sc_hd__dfxtp_1
X_13950_ _16099_/A vssd1 vssd1 vccd1 vccd1 _14333_/A sky130_fd_sc_hd__clkbuf_2
X_21059_ _21145_/A vssd1 vssd1 vccd1 vccd1 _21126_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25867_ _27154_/CLK _25867_/D vssd1 vssd1 vccd1 vccd1 _25867_/Q sky130_fd_sc_hd__dfxtp_1
X_13881_ _13920_/A vssd1 vssd1 vccd1 vccd1 _13891_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27606_ _27606_/CLK _27606_/D vssd1 vssd1 vccd1 vccd1 _27606_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _15620_/A vssd1 vssd1 vccd1 vccd1 _26171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24818_ _27638_/Q _24813_/X _24815_/Y _24817_/X vssd1 vssd1 vccd1 vccd1 _27638_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25798_ _25798_/A vssd1 vssd1 vccd1 vccd1 _27853_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27537_ _27608_/CLK _27537_/D vssd1 vssd1 vccd1 vccd1 _27537_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15551_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15608_/A sky130_fd_sc_hd__nor2_2
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24749_ _24940_/A vssd1 vssd1 vccd1 vccd1 _24759_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _26627_/Q _14496_/X _14492_/X _14501_/Y vssd1 vssd1 vccd1 vccd1 _26627_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _26955_/Q _26923_/Q _26891_/Q _26859_/Q _18244_/X _18269_/X vssd1 vssd1 vccd1
+ vccd1 _18270_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27468_ _27468_/CLK _27468_/D vssd1 vssd1 vccd1 vccd1 _27468_/Q sky130_fd_sc_hd__dfxtp_1
X_15482_ _13038_/X _26233_/Q _15490_/S vssd1 vssd1 vccd1 vccd1 _15483_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17221_ _17181_/X _17219_/X _17220_/X vssd1 vssd1 vccd1 vccd1 _17221_/X sky130_fd_sc_hd__a21bo_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14433_/A vssd1 vssd1 vccd1 vccd1 _15710_/A sky130_fd_sc_hd__buf_2
XFILLER_35_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26419_ _20769_/X _26419_/D vssd1 vssd1 vccd1 vccd1 _26419_/Q sky130_fd_sc_hd__dfxtp_1
X_27399_ _27401_/CLK _27399_/D vssd1 vssd1 vccd1 vccd1 _27399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17152_ _27206_/Q _17151_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17153_/A sky130_fd_sc_hd__mux2_1
X_14364_ _26669_/Q _14352_/X _14358_/X _14363_/Y vssd1 vssd1 vccd1 vccd1 _26669_/D
+ sky130_fd_sc_hd__a31o_1
Xinput15 la1_data_in[15] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_2
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 la1_data_in[25] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
Xinput37 la1_data_in[6] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_4
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 la1_oenb[16] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
X_16103_ _16369_/A vssd1 vssd1 vccd1 vccd1 _16360_/A sky130_fd_sc_hd__clkbuf_2
Xinput59 la1_oenb[26] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_4
X_13315_ _27003_/Q _13234_/X _13317_/S vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17083_ _17266_/A vssd1 vssd1 vccd1 vccd1 _17132_/S sky130_fd_sc_hd__clkbuf_2
X_14295_ _26694_/Q _14283_/X _14284_/X _14294_/Y vssd1 vssd1 vccd1 vccd1 _26694_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_143_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _16034_/A vssd1 vssd1 vccd1 vccd1 _16254_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_13246_ _15407_/A vssd1 vssd1 vccd1 vccd1 _14813_/B sky130_fd_sc_hd__buf_4
XFILLER_170_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13177_ _27345_/Q _13061_/A _13081_/A _27313_/Q _13176_/X vssd1 vssd1 vccd1 vccd1
+ _16169_/A sky130_fd_sc_hd__a221o_1
XFILLER_111_413 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17985_ _17830_/X _17984_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _17985_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19724_ _19710_/X _19711_/X _19712_/X _19713_/X _19714_/X _19715_/X vssd1 vssd1 vccd1
+ vccd1 _19725_/A sky130_fd_sc_hd__mux4_1
X_16936_ _27595_/Q _24208_/A _24207_/A _27594_/Q _16935_/X vssd1 vssd1 vccd1 vccd1
+ _16936_/X sky130_fd_sc_hd__o221a_1
XFILLER_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19655_ _19655_/A vssd1 vssd1 vccd1 vccd1 _19655_/X sky130_fd_sc_hd__clkbuf_1
X_16867_ _16867_/A _16867_/B vssd1 vssd1 vccd1 vccd1 _16867_/X sky130_fd_sc_hd__xor2_1
XFILLER_93_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18606_ _25564_/A vssd1 vssd1 vccd1 vccd1 _18606_/X sky130_fd_sc_hd__clkbuf_2
X_15818_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15827_/S sky130_fd_sc_hd__clkbuf_2
X_19586_ _19586_/A vssd1 vssd1 vccd1 vccd1 _19586_/X sky130_fd_sc_hd__clkbuf_1
X_16798_ _16798_/A _16798_/B vssd1 vssd1 vccd1 vccd1 _16798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18537_ _18468_/X _18532_/X _18536_/X _18412_/X vssd1 vssd1 vccd1 vccd1 _18546_/B
+ sky130_fd_sc_hd__a211o_1
X_15749_ _15749_/A _15758_/B vssd1 vssd1 vccd1 vccd1 _15749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18468_ _18468_/A vssd1 vssd1 vccd1 vccd1 _18468_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17419_ _17419_/A _17419_/B _17419_/C vssd1 vssd1 vccd1 vccd1 _23035_/C sky130_fd_sc_hd__nor3_2
X_18399_ _18399_/A vssd1 vssd1 vccd1 vccd1 _25966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20430_ _20500_/A vssd1 vssd1 vccd1 vccd1 _20430_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20361_ _25659_/A vssd1 vssd1 vccd1 vccd1 _20708_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22100_ _22100_/A vssd1 vssd1 vccd1 vccd1 _22100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23080_ _23080_/A vssd1 vssd1 vccd1 vccd1 _27084_/D sky130_fd_sc_hd__clkbuf_1
X_20292_ _20286_/X _20287_/X _20288_/X _20289_/X _20290_/X _20291_/X vssd1 vssd1 vccd1
+ vccd1 _20293_/A sky130_fd_sc_hd__mux4_1
X_22031_ _22016_/X _22018_/X _22020_/X _22022_/X _22023_/X _22024_/X vssd1 vssd1 vccd1
+ vccd1 _22032_/A sky130_fd_sc_hd__mux4_1
XFILLER_138_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26770_ _22006_/X _26770_/D vssd1 vssd1 vccd1 vccd1 _26770_/Q sky130_fd_sc_hd__dfxtp_1
X_23982_ _23943_/X _23980_/X _23981_/X _23958_/X vssd1 vssd1 vccd1 vccd1 _27294_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25721_ _25721_/A vssd1 vssd1 vccd1 vccd1 _25721_/X sky130_fd_sc_hd__clkbuf_1
X_22933_ _22923_/X _22924_/X _22925_/X _22926_/X _22927_/X _22928_/X vssd1 vssd1 vccd1
+ vccd1 _22934_/A sky130_fd_sc_hd__mux4_1
XFILLER_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25652_ _25652_/A vssd1 vssd1 vccd1 vccd1 _25652_/X sky130_fd_sc_hd__clkbuf_1
X_22864_ _22864_/A vssd1 vssd1 vccd1 vccd1 _22864_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24603_ _27661_/Q _24609_/B vssd1 vssd1 vccd1 vccd1 _24604_/A sky130_fd_sc_hd__and2_1
XFILLER_73_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21815_ _21809_/X _21810_/X _21811_/X _21812_/X _21813_/X _21814_/X vssd1 vssd1 vccd1
+ vccd1 _21816_/A sky130_fd_sc_hd__mux4_1
XFILLER_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25583_ _25583_/A vssd1 vssd1 vccd1 vccd1 _25583_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22795_ _22783_/X _22784_/X _22785_/X _22786_/X _22788_/X _22790_/X vssd1 vssd1 vccd1
+ vccd1 _22796_/A sky130_fd_sc_hd__mux4_1
XFILLER_184_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27322_ _27398_/CLK _27322_/D vssd1 vssd1 vccd1 vccd1 _27322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24534_ _27609_/Q vssd1 vssd1 vccd1 vccd1 _24534_/X sky130_fd_sc_hd__clkbuf_1
X_21746_ _21814_/A vssd1 vssd1 vccd1 vccd1 _21746_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27253_ _27776_/CLK _27253_/D vssd1 vssd1 vccd1 vccd1 _27253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24465_ _27630_/Q _24467_/B vssd1 vssd1 vccd1 vccd1 _24466_/A sky130_fd_sc_hd__and2_1
X_21677_ _21725_/A vssd1 vssd1 vccd1 vccd1 _21677_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26204_ _20027_/X _26204_/D vssd1 vssd1 vccd1 vccd1 _26204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23416_ _23416_/A _23416_/B _23507_/B vssd1 vssd1 vccd1 vccd1 _23485_/A sky130_fd_sc_hd__nor3b_1
X_20628_ _20617_/X _20619_/X _20621_/X _20623_/X _20624_/X _20625_/X vssd1 vssd1 vccd1
+ vccd1 _20629_/A sky130_fd_sc_hd__mux4_1
X_27184_ _27488_/CLK _27184_/D vssd1 vssd1 vccd1 vccd1 _27184_/Q sky130_fd_sc_hd__dfxtp_1
X_24396_ _24396_/A _24400_/B vssd1 vssd1 vccd1 vccd1 _24397_/A sky130_fd_sc_hd__and2_1
XFILLER_149_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26135_ _19787_/X _26135_/D vssd1 vssd1 vccd1 vccd1 _26135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20559_ _20559_/A vssd1 vssd1 vccd1 vccd1 _20559_/X sky130_fd_sc_hd__clkbuf_1
X_23347_ _24733_/A _27235_/Q _27248_/Q _24772_/A _23346_/Y vssd1 vssd1 vccd1 vccd1
+ _23360_/A sky130_fd_sc_hd__o221a_1
XFILLER_125_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13100_ _27058_/Q _13099_/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14080_ _14133_/A vssd1 vssd1 vccd1 vccd1 _14080_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26066_ _26069_/CLK _26066_/D vssd1 vssd1 vccd1 vccd1 _26066_/Q sky130_fd_sc_hd__dfxtp_1
X_23278_ _27725_/Q _23271_/Y _23277_/Y input57/X vssd1 vssd1 vccd1 vccd1 _23278_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13031_ _27368_/Q _27367_/Q vssd1 vssd1 vccd1 vccd1 _13231_/B sky130_fd_sc_hd__and2b_1
X_25017_ _25017_/A vssd1 vssd1 vccd1 vccd1 _27676_/D sky130_fd_sc_hd__clkbuf_1
X_22229_ _22261_/A vssd1 vssd1 vccd1 vccd1 _22229_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1075 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17770_ _25941_/Q _17769_/X _17770_/S vssd1 vssd1 vccd1 vccd1 _17771_/A sky130_fd_sc_hd__mux2_1
X_14982_ _26450_/Q _14974_/X _14976_/X _14981_/Y vssd1 vssd1 vccd1 vccd1 _26450_/D
+ sky130_fd_sc_hd__a31o_1
X_26968_ _22694_/X _26968_/D vssd1 vssd1 vccd1 vccd1 _26968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16721_ _16721_/A vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__inv_2
X_13933_ _14005_/A vssd1 vssd1 vccd1 vccd1 _13933_/X sky130_fd_sc_hd__clkbuf_2
X_25919_ _25985_/CLK _25919_/D vssd1 vssd1 vccd1 vccd1 _25919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26899_ _22450_/X _26899_/D vssd1 vssd1 vccd1 vccd1 _26899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19440_ _19524_/A _19440_/B vssd1 vssd1 vccd1 vccd1 _19440_/X sky130_fd_sc_hd__or2_1
X_16652_ _16652_/A _16652_/B vssd1 vssd1 vccd1 vccd1 _16654_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13864_ _14172_/A vssd1 vssd1 vccd1 vccd1 _13919_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15603_ _15603_/A vssd1 vssd1 vccd1 vccd1 _26179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19371_ _18929_/X _19370_/X _18932_/X vssd1 vssd1 vccd1 vccd1 _19371_/X sky130_fd_sc_hd__o21a_1
X_16583_ _16583_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _16588_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13795_ _13887_/A _13799_/B vssd1 vssd1 vccd1 vccd1 _13795_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18322_ _18322_/A vssd1 vssd1 vccd1 vccd1 _18322_/X sky130_fd_sc_hd__clkbuf_1
X_15534_ _13198_/X _26209_/Q _15534_/S vssd1 vssd1 vccd1 vccd1 _15535_/A sky130_fd_sc_hd__mux2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18253_ _18412_/A vssd1 vssd1 vccd1 vccd1 _18253_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _26240_/Q _13401_/X _15473_/S vssd1 vssd1 vccd1 vccd1 _15466_/A sky130_fd_sc_hd__mux2_1
XFILLER_187_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17204_ _27842_/Q _27146_/Q _25891_/Q _25859_/Q _17203_/X _17191_/X vssd1 vssd1 vccd1
+ vccd1 _17204_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14416_ _14532_/B vssd1 vssd1 vccd1 vccd1 _14416_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18184_ _18184_/A _18066_/X vssd1 vssd1 vccd1 vccd1 _18184_/X sky130_fd_sc_hd__or2b_1
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15396_ _15396_/A vssd1 vssd1 vccd1 vccd1 _26271_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1016 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17135_ _17120_/X _17134_/X _17098_/X vssd1 vssd1 vccd1 vccd1 _17135_/X sky130_fd_sc_hd__a21bo_1
X_14347_ _26676_/Q _14337_/X _14345_/X _14346_/Y vssd1 vssd1 vccd1 vccd1 _26676_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1049 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17066_ _17060_/X _17063_/X _17113_/S vssd1 vssd1 vccd1 vccd1 _17066_/X sky130_fd_sc_hd__mux2_1
X_14278_ _14304_/A vssd1 vssd1 vccd1 vccd1 _14289_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16017_ _27482_/Q _16017_/B vssd1 vssd1 vccd1 vccd1 _16017_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13229_ _27036_/Q _13228_/X _13229_/S vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__mux2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater402 _27357_/CLK vssd1 vssd1 vccd1 vccd1 _27338_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater413 _27311_/CLK vssd1 vssd1 vccd1 vccd1 _27386_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _17965_/X _17966_/X _18075_/S vssd1 vssd1 vccd1 vccd1 _17968_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_500 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater424 _26057_/CLK vssd1 vssd1 vccd1 vccd1 _27328_/CLK sky130_fd_sc_hd__clkbuf_1
X_19707_ _19707_/A vssd1 vssd1 vccd1 vccd1 _19707_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16919_ _16093_/X _16915_/Y _16918_/X vssd1 vssd1 vccd1 vccd1 _24261_/A sky130_fd_sc_hd__a21oi_2
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17899_ _18462_/A vssd1 vssd1 vccd1 vccd1 _17899_/X sky130_fd_sc_hd__buf_4
XFILLER_26_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19638_ _19638_/A vssd1 vssd1 vccd1 vccd1 _19638_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19569_ _19830_/A vssd1 vssd1 vccd1 vccd1 _19637_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21600_ _21648_/A vssd1 vssd1 vccd1 vccd1 _21600_/X sky130_fd_sc_hd__clkbuf_1
X_22580_ _22612_/A vssd1 vssd1 vccd1 vccd1 _22580_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21531_ _21563_/A vssd1 vssd1 vccd1 vccd1 _21531_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21462_ _21478_/A vssd1 vssd1 vccd1 vccd1 _21462_/X sky130_fd_sc_hd__clkbuf_1
X_24250_ _24250_/A _24250_/B vssd1 vssd1 vccd1 vccd1 _24251_/A sky130_fd_sc_hd__and2_1
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20413_ _20413_/A vssd1 vssd1 vccd1 vccd1 _20413_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23201_ _23201_/A vssd1 vssd1 vccd1 vccd1 _27137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21393_ _21651_/A vssd1 vssd1 vccd1 vccd1 _21463_/A sky130_fd_sc_hd__clkbuf_2
X_24181_ _24181_/A vssd1 vssd1 vccd1 vccd1 _27361_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20344_ _20334_/X _20335_/X _20336_/X _20337_/X _20339_/X _20341_/X vssd1 vssd1 vccd1
+ vccd1 _20345_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23132_ _27107_/Q _17705_/X _23132_/S vssd1 vssd1 vccd1 vccd1 _23133_/A sky130_fd_sc_hd__mux2_1
XFILLER_134_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27940_ _27940_/A _15942_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_23063_ _23063_/A vssd1 vssd1 vccd1 vccd1 _27076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20275_ _20323_/A vssd1 vssd1 vccd1 vccd1 _20275_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22014_ _22014_/A vssd1 vssd1 vccd1 vccd1 _22014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26822_ _22188_/X _26822_/D vssd1 vssd1 vccd1 vccd1 _26822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26753_ _21946_/X _26753_/D vssd1 vssd1 vccd1 vccd1 _26753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23965_ _27087_/Q _23954_/X _23955_/X _27119_/Q _23956_/X vssd1 vssd1 vccd1 vccd1
+ _23965_/X sky130_fd_sc_hd__a221o_1
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25704_ _25704_/A vssd1 vssd1 vccd1 vccd1 _25704_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22916_ _22916_/A vssd1 vssd1 vccd1 vccd1 _22916_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26684_ _21704_/X _26684_/D vssd1 vssd1 vccd1 vccd1 _26684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23896_ _23990_/A vssd1 vssd1 vccd1 vccd1 _23896_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25635_ _25635_/A vssd1 vssd1 vccd1 vccd1 _25635_/X sky130_fd_sc_hd__clkbuf_1
X_22847_ _22837_/X _22838_/X _22839_/X _22840_/X _22841_/X _22842_/X vssd1 vssd1 vccd1
+ vccd1 _22848_/A sky130_fd_sc_hd__mux4_1
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13639_/A vssd1 vssd1 vccd1 vccd1 _13580_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25566_ _27688_/Q vssd1 vssd1 vccd1 vccd1 _25566_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22778_ _22778_/A vssd1 vssd1 vccd1 vccd1 _22778_/X sky130_fd_sc_hd__clkbuf_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27305_ _27681_/CLK _27305_/D vssd1 vssd1 vccd1 vccd1 _27305_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24517_ _27607_/Q _24554_/B vssd1 vssd1 vccd1 vccd1 _24518_/A sky130_fd_sc_hd__and2_1
XFILLER_40_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21729_ _21721_/X _21722_/X _21723_/X _21724_/X _21725_/X _21726_/X vssd1 vssd1 vccd1
+ vccd1 _21730_/A sky130_fd_sc_hd__mux4_1
XFILLER_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25497_ _25592_/A vssd1 vssd1 vccd1 vccd1 _25497_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_427 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15250_ _14795_/X _26335_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15251_/A sky130_fd_sc_hd__mux2_1
X_27236_ _27236_/CLK _27236_/D vssd1 vssd1 vccd1 vccd1 _27236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24448_ _27622_/Q _24456_/B vssd1 vssd1 vccd1 vccd1 _24449_/A sky130_fd_sc_hd__and2_1
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14201_ _26728_/Q _14199_/X _14194_/X _14200_/Y vssd1 vssd1 vccd1 vccd1 _26728_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_184_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15181_ _15181_/A vssd1 vssd1 vccd1 vccd1 _26366_/D sky130_fd_sc_hd__clkbuf_1
X_27167_ _27225_/CLK _27167_/D vssd1 vssd1 vccd1 vccd1 _27167_/Q sky130_fd_sc_hd__dfxtp_1
X_24379_ _24379_/A vssd1 vssd1 vccd1 vccd1 _27471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14132_ _26753_/Q _14130_/X _14120_/X _14131_/Y vssd1 vssd1 vccd1 vccd1 _26753_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26118_ _19723_/X _26118_/D vssd1 vssd1 vccd1 vccd1 _26118_/Q sky130_fd_sc_hd__dfxtp_1
X_27098_ _27830_/CLK _27098_/D vssd1 vssd1 vccd1 vccd1 _27098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _14079_/A vssd1 vssd1 vccd1 vccd1 _14147_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18940_ _26686_/Q _26654_/Q _26622_/Q _26590_/Q _18847_/X _18939_/X vssd1 vssd1 vccd1
+ vccd1 _18940_/X sky130_fd_sc_hd__mux4_2
X_26049_ _26049_/CLK _26049_/D vssd1 vssd1 vccd1 vccd1 _26049_/Q sky130_fd_sc_hd__dfxtp_1
X_13014_ _13014_/A vssd1 vssd1 vccd1 vccd1 _27793_/D sky130_fd_sc_hd__clkbuf_1
X_18871_ _26812_/Q _26780_/Q _26748_/Q _26716_/Q _18870_/X _18770_/X vssd1 vssd1 vccd1
+ vccd1 _18872_/B sky130_fd_sc_hd__mux4_1
XFILLER_67_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17822_ _17898_/A vssd1 vssd1 vccd1 vccd1 _18403_/A sky130_fd_sc_hd__buf_2
XFILLER_79_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17753_ _27432_/Q vssd1 vssd1 vccd1 vccd1 _17753_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14965_ _26456_/Q _14957_/X _14960_/X _14964_/Y vssd1 vssd1 vccd1 vccd1 _26456_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13916_ _26820_/Q _13906_/X _13912_/X _13915_/Y vssd1 vssd1 vccd1 vccd1 _26820_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16704_ _16076_/A _16744_/A _16372_/A _16084_/A vssd1 vssd1 vccd1 vccd1 _16704_/X
+ sky130_fd_sc_hd__a31o_1
X_17684_ _25914_/Q _17683_/X _17690_/S vssd1 vssd1 vccd1 vccd1 _17685_/A sky130_fd_sc_hd__mux2_1
X_14896_ _14724_/X _26485_/Q _14896_/S vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__mux2_1
X_16635_ _16619_/X _16631_/Y _16634_/X _16626_/X vssd1 vssd1 vccd1 vccd1 _24247_/A
+ sky130_fd_sc_hd__a22o_1
X_19423_ _26546_/Q _26514_/Q _26482_/Q _27058_/Q _19401_/X _19287_/X vssd1 vssd1 vccd1
+ vccd1 _19423_/X sky130_fd_sc_hd__mux4_1
X_13847_ _13940_/A _13847_/B vssd1 vssd1 vccd1 vccd1 _13847_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16566_ _16301_/B _16301_/C _16576_/A vssd1 vssd1 vccd1 vccd1 _16567_/B sky130_fd_sc_hd__o21ai_1
XFILLER_16_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19354_ _19488_/A vssd1 vssd1 vccd1 vccd1 _19354_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13778_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13778_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15517_ _13150_/X _26217_/Q _15523_/S vssd1 vssd1 vccd1 vccd1 _15518_/A sky130_fd_sc_hd__mux2_1
X_18305_ _18305_/A vssd1 vssd1 vccd1 vccd1 _18305_/X sky130_fd_sc_hd__buf_2
XFILLER_188_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19285_ _19191_/X _19284_/X _19194_/X vssd1 vssd1 vccd1 vccd1 _19285_/X sky130_fd_sc_hd__o21a_1
XFILLER_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16497_ _16697_/A _16497_/B vssd1 vssd1 vccd1 vccd1 _16499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_176_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ _18395_/A vssd1 vssd1 vccd1 vccd1 _18331_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15448_ _15448_/A vssd1 vssd1 vccd1 vccd1 _26248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ _18165_/X _18166_/X _18216_/S vssd1 vssd1 vccd1 vccd1 _18167_/X sky130_fd_sc_hd__mux2_2
XFILLER_117_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ _14772_/X _26278_/Q _15379_/S vssd1 vssd1 vccd1 vccd1 _15380_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17118_ _25921_/Q _25987_/Q _17132_/S vssd1 vssd1 vccd1 vccd1 _17119_/B sky130_fd_sc_hd__mux2_1
XFILLER_156_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18098_ _18098_/A vssd1 vssd1 vccd1 vccd1 _25953_/D sky130_fd_sc_hd__clkbuf_1
X_17049_ _27198_/Q _17048_/X _17067_/S vssd1 vssd1 vccd1 vccd1 _17050_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20060_ _20076_/A vssd1 vssd1 vccd1 vccd1 _20060_/X sky130_fd_sc_hd__clkbuf_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater210 _25913_/CLK vssd1 vssd1 vccd1 vccd1 _27417_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater221 _27404_/CLK vssd1 vssd1 vccd1 vccd1 _27401_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater232 _27602_/CLK vssd1 vssd1 vccd1 vccd1 _27601_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater243 _27623_/CLK vssd1 vssd1 vccd1 vccd1 _27625_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater254 _27617_/CLK vssd1 vssd1 vccd1 vccd1 _27621_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater265 _27593_/CLK vssd1 vssd1 vccd1 vccd1 _27185_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater276 _27539_/CLK vssd1 vssd1 vccd1 vccd1 _27541_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23750_ _25912_/Q _25978_/Q _25811_/Q _26010_/Q _23747_/X _23749_/X vssd1 vssd1 vccd1
+ vccd1 _23750_/X sky130_fd_sc_hd__mux4_1
Xrepeater287 _27477_/CLK vssd1 vssd1 vccd1 vccd1 _27372_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _20962_/A vssd1 vssd1 vccd1 vccd1 _20962_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater298 _27236_/CLK vssd1 vssd1 vccd1 vccd1 _27264_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22701_ _22959_/A vssd1 vssd1 vccd1 vccd1 _22771_/A sky130_fd_sc_hd__buf_2
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23681_ _27766_/Q _27246_/Q _23683_/S vssd1 vssd1 vccd1 vccd1 _23682_/A sky130_fd_sc_hd__mux2_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20893_ _20941_/A vssd1 vssd1 vccd1 vccd1 _20893_/X sky130_fd_sc_hd__clkbuf_2
X_25420_ _27748_/Q input60/X _25424_/S vssd1 vssd1 vccd1 vccd1 _25421_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22632_ _22698_/A vssd1 vssd1 vccd1 vccd1 _22632_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25351_ _25356_/A _25351_/B vssd1 vssd1 vccd1 vccd1 _25351_/Y sky130_fd_sc_hd__nand2_1
X_22563_ _22611_/A vssd1 vssd1 vccd1 vccd1 _22563_/X sky130_fd_sc_hd__clkbuf_1
X_24302_ _24302_/A _24302_/B vssd1 vssd1 vccd1 vccd1 _27432_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21514_ _21562_/A vssd1 vssd1 vccd1 vccd1 _21514_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25282_ _25282_/A _25282_/B vssd1 vssd1 vccd1 vccd1 _25283_/B sky130_fd_sc_hd__xnor2_1
X_22494_ _22494_/A vssd1 vssd1 vccd1 vccd1 _22494_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27021_ _22880_/X _27021_/D vssd1 vssd1 vccd1 vccd1 _27021_/Q sky130_fd_sc_hd__dfxtp_1
X_24233_ _24233_/A _24233_/B vssd1 vssd1 vccd1 vccd1 _24234_/A sky130_fd_sc_hd__and2_1
X_21445_ _21477_/A vssd1 vssd1 vccd1 vccd1 _21445_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21376_ _21392_/A vssd1 vssd1 vccd1 vccd1 _21376_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24164_ _24175_/A vssd1 vssd1 vccd1 vccd1 _24173_/B sky130_fd_sc_hd__clkbuf_1
X_20327_ _20327_/A vssd1 vssd1 vccd1 vccd1 _20327_/X sky130_fd_sc_hd__clkbuf_1
X_23115_ _27099_/Q _17680_/X _23121_/S vssd1 vssd1 vccd1 vccd1 _23116_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24095_ _27396_/Q _24095_/B vssd1 vssd1 vccd1 vccd1 _24096_/A sky130_fd_sc_hd__and2_1
XFILLER_162_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20258_ _20248_/X _20249_/X _20250_/X _20251_/X _20253_/X _20255_/X vssd1 vssd1 vccd1
+ vccd1 _20259_/A sky130_fd_sc_hd__mux4_1
X_27923_ _27923_/A _15964_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
X_23046_ _27069_/Q _17686_/X _23048_/S vssd1 vssd1 vccd1 vccd1 _23047_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27854_ _27854_/CLK _27854_/D vssd1 vssd1 vccd1 vccd1 _27854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20189_ _20237_/A vssd1 vssd1 vccd1 vccd1 _20189_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26805_ _22132_/X _26805_/D vssd1 vssd1 vccd1 vccd1 _26805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27785_ _27787_/CLK _27785_/D vssd1 vssd1 vccd1 vccd1 _27785_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24997_ _25103_/S vssd1 vssd1 vccd1 vccd1 _25031_/S sky130_fd_sc_hd__buf_2
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26736_ _21888_/X _26736_/D vssd1 vssd1 vccd1 vccd1 _26736_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14750_/A vssd1 vssd1 vccd1 vccd1 _14750_/X sky130_fd_sc_hd__buf_2
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23948_ _27787_/Q vssd1 vssd1 vccd1 vccd1 _23985_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13882_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13701_/Y sky130_fd_sc_hd__nor2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26667_ _21642_/X _26667_/D vssd1 vssd1 vccd1 vccd1 _26667_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _26565_/Q _14671_/X _14679_/X _14680_/Y vssd1 vssd1 vccd1 vccd1 _26565_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23879_ _27078_/Q _23860_/X _23861_/X _27110_/Q _23862_/X vssd1 vssd1 vccd1 vccd1
+ _23879_/X sky130_fd_sc_hd__a221o_1
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16420_ _16420_/A _16508_/B vssd1 vssd1 vccd1 vccd1 _16420_/Y sky130_fd_sc_hd__nor2_1
X_13632_ _13902_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13632_/Y sky130_fd_sc_hd__nor2_1
X_25618_ _25618_/A _25618_/B vssd1 vssd1 vccd1 vccd1 _27788_/D sky130_fd_sc_hd__nor2_1
XFILLER_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26598_ _21404_/X _26598_/D vssd1 vssd1 vccd1 vccd1 _26598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16351_ _16754_/A _16351_/B vssd1 vssd1 vccd1 vccd1 _16857_/A sky130_fd_sc_hd__and2_1
X_25549_ _25530_/X _25261_/B _25548_/X _25543_/X vssd1 vssd1 vccd1 vccd1 _25549_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ _27339_/Q _13529_/X _13530_/X _27307_/Q _13213_/X vssd1 vssd1 vccd1 vccd1
+ _14518_/A sky130_fd_sc_hd__a221oi_4
XFILLER_157_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15302_ _26312_/Q _13376_/X _15306_/S vssd1 vssd1 vccd1 vccd1 _15303_/A sky130_fd_sc_hd__mux2_1
XFILLER_201_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19070_ _19482_/A vssd1 vssd1 vccd1 vccd1 _19070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16282_ _26062_/Q vssd1 vssd1 vccd1 vccd1 _16282_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13494_ _13891_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18021_ _26272_/Q _26240_/Q _26208_/Q _26176_/Q _17873_/X _17937_/X vssd1 vssd1 vccd1
+ vccd1 _18021_/X sky130_fd_sc_hd__mux4_1
X_27219_ _27219_/CLK _27219_/D vssd1 vssd1 vccd1 vccd1 _27219_/Q sky130_fd_sc_hd__dfxtp_1
X_15233_ _15233_/A vssd1 vssd1 vccd1 vccd1 _26343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15164_ _15175_/A vssd1 vssd1 vccd1 vccd1 _15173_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_197_1092 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14115_ _14381_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15095_ _14779_/X _26404_/Q _15101_/S vssd1 vssd1 vccd1 vccd1 _15096_/A sky130_fd_sc_hd__mux2_1
X_19972_ _19988_/A vssd1 vssd1 vccd1 vccd1 _19972_/X sky130_fd_sc_hd__clkbuf_1
X_14046_ _14518_/A vssd1 vssd1 vccd1 vccd1 _14403_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18923_ _18923_/A vssd1 vssd1 vccd1 vccd1 _18923_/X sky130_fd_sc_hd__buf_4
XFILLER_68_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18854_ _19324_/A vssd1 vssd1 vccd1 vccd1 _18854_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17805_ _18012_/A vssd1 vssd1 vccd1 vccd1 _17805_/X sky130_fd_sc_hd__buf_4
X_15997_ _27479_/Q _27370_/Q vssd1 vssd1 vccd1 vccd1 _16001_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18785_ _18932_/A vssd1 vssd1 vccd1 vccd1 _18785_/X sky130_fd_sc_hd__buf_2
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17736_ _17736_/A vssd1 vssd1 vccd1 vccd1 _25930_/D sky130_fd_sc_hd__clkbuf_1
X_14948_ _14948_/A vssd1 vssd1 vccd1 vccd1 _26462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17667_ _17517_/X _25904_/Q _17667_/S vssd1 vssd1 vccd1 vccd1 _17668_/A sky130_fd_sc_hd__mux2_1
X_14879_ _26492_/Q _13414_/X _14879_/S vssd1 vssd1 vccd1 vccd1 _14880_/A sky130_fd_sc_hd__mux2_1
X_19406_ _19406_/A vssd1 vssd1 vccd1 vccd1 _26065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16618_ _16660_/A _16618_/B vssd1 vssd1 vccd1 vccd1 _16618_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17598_ _17598_/A vssd1 vssd1 vccd1 vccd1 _25873_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16549_ _16662_/A _16911_/A vssd1 vssd1 vccd1 vccd1 _16549_/X sky130_fd_sc_hd__and2_1
X_19337_ _19337_/A vssd1 vssd1 vccd1 vccd1 _26062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19268_ _19362_/A _19268_/B _19268_/C vssd1 vssd1 vccd1 vccd1 _19269_/A sky130_fd_sc_hd__and3_1
XFILLER_148_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18219_/A vssd1 vssd1 vccd1 vccd1 _25958_/D sky130_fd_sc_hd__clkbuf_1
X_19199_ _19196_/X _19197_/X _19334_/S vssd1 vssd1 vccd1 vccd1 _19199_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21230_ _21579_/A vssd1 vssd1 vccd1 vccd1 _21301_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21161_ _21144_/X _21146_/X _21148_/X _21150_/X _21151_/X _21152_/X vssd1 vssd1 vccd1
+ vccd1 _21162_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20112_ _20095_/X _20097_/X _20099_/X _20101_/X _20102_/X _20103_/X vssd1 vssd1 vccd1
+ vccd1 _20113_/A sky130_fd_sc_hd__mux4_1
X_21092_ _21092_/A vssd1 vssd1 vccd1 vccd1 _21092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20043_ _20043_/A vssd1 vssd1 vccd1 vccd1 _20043_/X sky130_fd_sc_hd__clkbuf_1
X_24920_ _24937_/A _24920_/B vssd1 vssd1 vccd1 vccd1 _24920_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24851_ _27760_/Q _27759_/Q _24851_/C vssd1 vssd1 vccd1 vccd1 _24857_/B sky130_fd_sc_hd__and3_1
XFILLER_74_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23802_ _23991_/A vssd1 vssd1 vccd1 vccd1 _23802_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27570_ _27577_/CLK _27570_/D vssd1 vssd1 vccd1 vccd1 _27570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24782_ _24782_/A _24786_/B vssd1 vssd1 vccd1 vccd1 _24782_/Y sky130_fd_sc_hd__nand2_1
X_21994_ _21994_/A vssd1 vssd1 vccd1 vccd1 _21994_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _22613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26521_ _21136_/X _26521_/D vssd1 vssd1 vccd1 vccd1 _26521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _22543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_23733_ _23733_/A vssd1 vssd1 vccd1 vccd1 _27268_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_129 _24925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20945_ _20937_/X _20938_/X _20939_/X _20940_/X _20941_/X _20942_/X vssd1 vssd1 vccd1
+ vccd1 _20946_/A sky130_fd_sc_hd__mux4_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26452_ _20900_/X _26452_/D vssd1 vssd1 vccd1 vccd1 _26452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23664_ _24844_/A _27238_/Q _23672_/S vssd1 vssd1 vccd1 vccd1 _23665_/A sky130_fd_sc_hd__mux2_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20876_ _20876_/A vssd1 vssd1 vccd1 vccd1 _20876_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25403_ _25403_/A vssd1 vssd1 vccd1 vccd1 _27740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_197_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22615_ _22685_/A vssd1 vssd1 vccd1 vccd1 _22615_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26383_ _20649_/X _26383_/D vssd1 vssd1 vccd1 vccd1 _26383_/Q sky130_fd_sc_hd__dfxtp_1
X_23595_ _25580_/A _27219_/Q _23595_/S vssd1 vssd1 vccd1 vccd1 _23596_/B sky130_fd_sc_hd__mux2_1
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25334_ _25331_/Y _25332_/X _25329_/X _25330_/Y _25319_/C vssd1 vssd1 vccd1 vccd1
+ _25335_/B sky130_fd_sc_hd__o2111ai_1
XFILLER_195_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22546_ _22546_/A vssd1 vssd1 vccd1 vccd1 _22893_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25265_ _25265_/A _25265_/B vssd1 vssd1 vccd1 vccd1 _25265_/Y sky130_fd_sc_hd__nor2_1
X_22477_ _22471_/X _22472_/X _22473_/X _22474_/X _22475_/X _22476_/X vssd1 vssd1 vccd1
+ vccd1 _22478_/A sky130_fd_sc_hd__mux4_1
XFILLER_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27004_ _22820_/X _27004_/D vssd1 vssd1 vccd1 vccd1 _27004_/Q sky130_fd_sc_hd__dfxtp_1
X_24216_ _24216_/A vssd1 vssd1 vccd1 vccd1 _27376_/D sky130_fd_sc_hd__clkbuf_1
X_21428_ _21476_/A vssd1 vssd1 vccd1 vccd1 _21428_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25196_ _27530_/Q _27498_/Q vssd1 vssd1 vccd1 vccd1 _25197_/B sky130_fd_sc_hd__or2_1
XFILLER_146_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_677 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24147_ _27451_/Q _24151_/B vssd1 vssd1 vccd1 vccd1 _24148_/A sky130_fd_sc_hd__and2_1
X_21359_ _21391_/A vssd1 vssd1 vccd1 vccd1 _21359_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24078_ _27388_/Q _24084_/B vssd1 vssd1 vccd1 vccd1 _24079_/A sky130_fd_sc_hd__and2_1
XFILLER_122_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15920_ _15924_/A vssd1 vssd1 vccd1 vccd1 _15920_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23029_ _23029_/A vssd1 vssd1 vccd1 vccd1 _23029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1026 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15851_ _13234_/X _26075_/Q _15853_/S vssd1 vssd1 vccd1 vccd1 _15852_/A sky130_fd_sc_hd__mux2_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27837_ _27837_/CLK _27837_/D vssd1 vssd1 vccd1 vccd1 _27837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14801_/X _26525_/Q _14805_/S vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__mux2_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18570_ _26713_/Q _26681_/Q _26649_/Q _26617_/Q _18345_/X _18012_/A vssd1 vssd1 vccd1
+ vccd1 _18571_/A sky130_fd_sc_hd__mux4_1
X_15782_ _26106_/Q _15774_/X _15703_/B _15781_/Y vssd1 vssd1 vccd1 vccd1 _26106_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_188_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _27801_/Q _12998_/B vssd1 vssd1 vccd1 vccd1 _12995_/A sky130_fd_sc_hd__and2_1
X_27768_ _27768_/CLK _27768_/D vssd1 vssd1 vccd1 vccd1 _27768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ _17520_/X _25841_/Q _17524_/S vssd1 vssd1 vccd1 vccd1 _17522_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _14733_/A vssd1 vssd1 vccd1 vccd1 _26547_/D sky130_fd_sc_hd__clkbuf_1
X_26719_ _21824_/X _26719_/D vssd1 vssd1 vccd1 vccd1 _26719_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27984__450 vssd1 vssd1 vccd1 vccd1 _27984__450/HI _27984_/A sky130_fd_sc_hd__conb_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27699_ _27699_/CLK _27699_/D vssd1 vssd1 vccd1 vccd1 _27699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17452_ _17452_/A vssd1 vssd1 vccd1 vccd1 _25819_/D sky130_fd_sc_hd__clkbuf_1
X_14664_ _15738_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14664_/Y sky130_fd_sc_hd__nor2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _27385_/Q _16557_/B vssd1 vssd1 vccd1 vccd1 _16403_/Y sky130_fd_sc_hd__nand2_1
X_13615_ _26928_/Q _13613_/X _13603_/X _13614_/Y vssd1 vssd1 vccd1 vccd1 _26928_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_189_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17383_ _16992_/X _17382_/X _17342_/X vssd1 vssd1 vccd1 vccd1 _17383_/X sky130_fd_sc_hd__a21bo_1
X_14595_ _15756_/A _14597_/B vssd1 vssd1 vccd1 vccd1 _14595_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19122_ _26149_/Q _26085_/Q _27013_/Q _26981_/Q _19049_/X _19070_/X vssd1 vssd1 vccd1
+ vccd1 _19123_/B sky130_fd_sc_hd__mux4_1
X_16334_ _14804_/A _16501_/A _16412_/A _25946_/Q _16333_/Y vssd1 vssd1 vccd1 vccd1
+ _16756_/B sky130_fd_sc_hd__a221o_1
X_13546_ _13546_/A vssd1 vssd1 vccd1 vccd1 _13565_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19053_ _18954_/X _19052_/X _18958_/X vssd1 vssd1 vccd1 vccd1 _19053_/X sky130_fd_sc_hd__o21a_1
X_16265_ _16263_/Y _16119_/A _16277_/B _16495_/A _16264_/Y vssd1 vssd1 vccd1 vccd1
+ _24293_/A sky130_fd_sc_hd__o221a_1
X_13477_ _26961_/Q _13464_/X _13457_/X _13476_/Y vssd1 vssd1 vccd1 vccd1 _26961_/D
+ sky130_fd_sc_hd__a31o_1
X_15216_ _15216_/A vssd1 vssd1 vccd1 vccd1 _26351_/D sky130_fd_sc_hd__clkbuf_1
X_18004_ _18458_/A vssd1 vssd1 vccd1 vccd1 _18004_/X sky130_fd_sc_hd__buf_4
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16196_ _17410_/A _16224_/B vssd1 vssd1 vccd1 vccd1 _16196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ _26381_/Q _13360_/X _15151_/S vssd1 vssd1 vccd1 vccd1 _15148_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19955_ _19955_/A vssd1 vssd1 vccd1 vccd1 _19955_/X sky130_fd_sc_hd__clkbuf_1
X_15078_ _15078_/A vssd1 vssd1 vccd1 vccd1 _26412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27952__438 vssd1 vssd1 vccd1 vccd1 _27952__438/HI _27952_/A sky130_fd_sc_hd__conb_1
X_14029_ _14390_/A _14029_/B vssd1 vssd1 vccd1 vccd1 _14029_/Y sky130_fd_sc_hd__nor2_1
X_18906_ _19431_/A vssd1 vssd1 vccd1 vccd1 _19501_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19886_ _19886_/A vssd1 vssd1 vccd1 vccd1 _19886_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18837_ _19290_/A vssd1 vssd1 vccd1 vccd1 _18837_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18768_ _27599_/Q vssd1 vssd1 vccd1 vccd1 _19460_/A sky130_fd_sc_hd__buf_2
X_17719_ _25925_/Q _17718_/X _17722_/S vssd1 vssd1 vccd1 vccd1 _17720_/A sky130_fd_sc_hd__mux2_1
X_18699_ _18699_/A vssd1 vssd1 vccd1 vccd1 _26012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20730_ _20722_/X _20723_/X _20724_/X _20725_/X _20726_/X _20727_/X vssd1 vssd1 vccd1
+ vccd1 _20731_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20661_ _20661_/A vssd1 vssd1 vccd1 vccd1 _20661_/X sky130_fd_sc_hd__clkbuf_1
X_22400_ _22400_/A vssd1 vssd1 vccd1 vccd1 _22400_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20592_ _20582_/X _20583_/X _20584_/X _20585_/X _20586_/X _20587_/X vssd1 vssd1 vccd1
+ vccd1 _20593_/A sky130_fd_sc_hd__mux4_2
X_23380_ _24825_/A _27234_/Q _27245_/Q _24765_/A vssd1 vssd1 vccd1 vccd1 _23380_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22331_ _22347_/A vssd1 vssd1 vccd1 vccd1 _22331_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25050_ _25050_/A vssd1 vssd1 vccd1 vccd1 _27680_/D sky130_fd_sc_hd__clkbuf_1
X_22262_ _22262_/A vssd1 vssd1 vccd1 vccd1 _22262_/X sky130_fd_sc_hd__clkbuf_1
X_24001_ _24001_/A vssd1 vssd1 vccd1 vccd1 _24001_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21213_ _21213_/A vssd1 vssd1 vccd1 vccd1 _21213_/X sky130_fd_sc_hd__clkbuf_1
X_22193_ _22451_/A vssd1 vssd1 vccd1 vccd1 _22261_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_400 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21144_ _21211_/A vssd1 vssd1 vccd1 vccd1 _21144_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21075_ _21058_/X _21060_/X _21062_/X _21064_/X _21065_/X _21066_/X vssd1 vssd1 vccd1
+ vccd1 _21076_/A sky130_fd_sc_hd__mux4_1
X_25952_ _25953_/CLK _25952_/D vssd1 vssd1 vccd1 vccd1 _25952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_499 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24903_ _24910_/C _24903_/B vssd1 vssd1 vccd1 vccd1 _24904_/B sky130_fd_sc_hd__or2_1
X_20026_ _20009_/X _20011_/X _20013_/X _20015_/X _20016_/X _20017_/X vssd1 vssd1 vccd1
+ vccd1 _20027_/A sky130_fd_sc_hd__mux4_1
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25883_ _25884_/CLK _25883_/D vssd1 vssd1 vccd1 vccd1 _25883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27622_ _27700_/CLK _27622_/D vssd1 vssd1 vccd1 vccd1 _27622_/Q sky130_fd_sc_hd__dfxtp_1
X_24834_ _24861_/A vssd1 vssd1 vccd1 vccd1 _24834_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27553_ _27555_/CLK _27553_/D vssd1 vssd1 vccd1 vccd1 _27553_/Q sky130_fd_sc_hd__dfxtp_1
X_24765_ _24765_/A _24772_/B vssd1 vssd1 vccd1 vccd1 _24765_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ _21965_/X _21966_/X _21967_/X _21968_/X _21969_/X _21970_/X vssd1 vssd1 vccd1
+ vccd1 _21978_/A sky130_fd_sc_hd__mux4_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26504_ _21076_/X _26504_/D vssd1 vssd1 vccd1 vccd1 _26504_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23716_ _24960_/A _27262_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23717_/A sky130_fd_sc_hd__mux2_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20928_ _20928_/A vssd1 vssd1 vccd1 vccd1 _20928_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27484_ _27484_/CLK _27484_/D vssd1 vssd1 vccd1 vccd1 _27484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24696_ _27180_/Q _24698_/B vssd1 vssd1 vccd1 vccd1 _24696_/X sky130_fd_sc_hd__or2_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26435_ _20839_/X _26435_/D vssd1 vssd1 vccd1 vccd1 _26435_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23647_ _23643_/X _23638_/X _24987_/S vssd1 vssd1 vccd1 vccd1 _23649_/A sky130_fd_sc_hd__a21oi_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20859_ _20859_/A vssd1 vssd1 vccd1 vccd1 _20859_/X sky130_fd_sc_hd__clkbuf_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ _13400_/A vssd1 vssd1 vccd1 vccd1 _26977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_186_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14380_ _14393_/A vssd1 vssd1 vccd1 vccd1 _14390_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_26366_ _20591_/X _26366_/D vssd1 vssd1 vccd1 vccd1 _26366_/Q sky130_fd_sc_hd__dfxtp_1
X_23578_ _23578_/A vssd1 vssd1 vccd1 vccd1 _27214_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25317_ _25323_/A _27513_/Q vssd1 vssd1 vccd1 vccd1 _25328_/A sky130_fd_sc_hd__xnor2_1
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13331_ _14721_/A vssd1 vssd1 vccd1 vccd1 _13331_/X sky130_fd_sc_hd__buf_2
XFILLER_167_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22529_ _22519_/X _22520_/X _22521_/X _22522_/X _22524_/X _22526_/X vssd1 vssd1 vccd1
+ vccd1 _22530_/A sky130_fd_sc_hd__mux4_1
XFILLER_127_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26297_ _20347_/X _26297_/D vssd1 vssd1 vccd1 vccd1 _26297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16050_ _16047_/Y _27370_/Q _16048_/X _16049_/Y _27369_/Q vssd1 vssd1 vccd1 vccd1
+ _16066_/C sky130_fd_sc_hd__o221a_1
XFILLER_157_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25248_ _27537_/Q _27505_/Q vssd1 vssd1 vccd1 vccd1 _25267_/A sky130_fd_sc_hd__nand2_1
X_13262_ _13262_/A vssd1 vssd1 vccd1 vccd1 _27028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15001_ _25106_/A vssd1 vssd1 vccd1 vccd1 _15705_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25179_ _25190_/A _25179_/B vssd1 vssd1 vccd1 vccd1 _25181_/A sky130_fd_sc_hd__nand2_1
X_13193_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13193_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19740_ _19726_/X _19727_/X _19728_/X _19729_/X _19731_/X _19733_/X vssd1 vssd1 vccd1
+ vccd1 _19741_/A sky130_fd_sc_hd__mux4_1
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16952_ _27584_/Q vssd1 vssd1 vccd1 vccd1 _24633_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15903_ _15906_/A vssd1 vssd1 vccd1 vccd1 _15903_/Y sky130_fd_sc_hd__inv_2
X_19671_ _19671_/A vssd1 vssd1 vccd1 vccd1 _19671_/X sky130_fd_sc_hd__clkbuf_1
X_16883_ _16877_/X _16879_/X _16880_/Y _16882_/X vssd1 vssd1 vccd1 vccd1 _24262_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18622_ _25978_/Q _17673_/X _18630_/S vssd1 vssd1 vccd1 vccd1 _18623_/A sky130_fd_sc_hd__mux2_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _13184_/X _26083_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15835_/A sky130_fd_sc_hd__mux2_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18553_/A _18474_/X vssd1 vssd1 vccd1 vccd1 _18553_/X sky130_fd_sc_hd__or2b_1
XFILLER_79_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _26113_/Q _15760_/X _15753_/X _15764_/Y vssd1 vssd1 vccd1 vccd1 _26113_/D
+ sky130_fd_sc_hd__a31o_1
X_12977_ _12977_/A vssd1 vssd1 vccd1 vccd1 _27809_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _27433_/Q vssd1 vssd1 vccd1 vccd1 _17504_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14716_ _14715_/X _26552_/Q _14725_/S vssd1 vssd1 vccd1 vccd1 _14717_/A sky130_fd_sc_hd__mux2_1
X_15696_ _15712_/A vssd1 vssd1 vccd1 vccd1 _15781_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18484_ _18437_/X _18482_/X _18483_/X vssd1 vssd1 vccd1 vccd1 _18484_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _26578_/Q _14645_/X _14640_/X _14646_/Y vssd1 vssd1 vccd1 vccd1 _26578_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17435_ _17434_/X _25814_/Q _17438_/S vssd1 vssd1 vccd1 vccd1 _17436_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_18 _25992_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14578_ _26603_/Q _14576_/X _14566_/X _14577_/Y vssd1 vssd1 vccd1 vccd1 _26603_/D
+ sky130_fd_sc_hd__a31o_1
X_17366_ _17364_/X _17365_/X _17386_/S vssd1 vssd1 vccd1 vccd1 _17366_/X sky130_fd_sc_hd__mux2_2
XANTENNA_29 _27836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19105_ _19220_/A vssd1 vssd1 vccd1 vccd1 _19105_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16317_ _16792_/B vssd1 vssd1 vccd1 vccd1 _16598_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13529_ _13529_/A vssd1 vssd1 vccd1 vccd1 _13529_/X sky130_fd_sc_hd__buf_4
X_17297_ _27218_/Q _17296_/X _17311_/S vssd1 vssd1 vccd1 vccd1 _17298_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19036_ _19027_/X _19030_/X _19034_/X _19035_/X _18987_/X vssd1 vssd1 vccd1 vccd1
+ _19037_/C sky130_fd_sc_hd__a221o_1
X_16248_ _16728_/A _16460_/B vssd1 vssd1 vccd1 vccd1 _16256_/C sky130_fd_sc_hd__or2_1
XFILLER_161_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16179_ _16172_/X _16173_/X _16176_/Y _16177_/X _16178_/X vssd1 vssd1 vccd1 vccd1
+ _16345_/A sky130_fd_sc_hd__o41a_1
XFILLER_99_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19938_ _19918_/X _19921_/X _19924_/X _19927_/X _19928_/X _19929_/X vssd1 vssd1 vccd1
+ vccd1 _19939_/A sky130_fd_sc_hd__mux4_1
X_19869_ _19901_/A vssd1 vssd1 vccd1 vccd1 _19869_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21900_ _21900_/A vssd1 vssd1 vccd1 vccd1 _21900_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22880_ _22880_/A vssd1 vssd1 vccd1 vccd1 _22880_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21831_ _22089_/A vssd1 vssd1 vccd1 vccd1 _21900_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24550_ _24550_/A vssd1 vssd1 vccd1 vccd1 _27537_/D sky130_fd_sc_hd__clkbuf_1
X_21762_ _21827_/A vssd1 vssd1 vccd1 vccd1 _21762_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23501_ input33/X _23429_/A _23500_/X _23498_/X vssd1 vssd1 vccd1 vccd1 _27193_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20713_ _20713_/A vssd1 vssd1 vccd1 vccd1 _20713_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24481_ _27637_/Q _24509_/B vssd1 vssd1 vccd1 vccd1 _24482_/A sky130_fd_sc_hd__and2_1
X_21693_ _21725_/A vssd1 vssd1 vccd1 vccd1 _21693_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26220_ _20085_/X _26220_/D vssd1 vssd1 vccd1 vccd1 _26220_/Q sky130_fd_sc_hd__dfxtp_1
X_23432_ _23500_/B vssd1 vssd1 vccd1 vccd1 _23443_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_20644_ _20636_/X _20637_/X _20638_/X _20639_/X _20640_/X _20641_/X vssd1 vssd1 vccd1
+ vccd1 _20645_/A sky130_fd_sc_hd__mux4_1
XFILLER_20_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26151_ _19843_/X _26151_/D vssd1 vssd1 vccd1 vccd1 _26151_/Q sky130_fd_sc_hd__dfxtp_1
X_23363_ _27259_/Q vssd1 vssd1 vccd1 vccd1 _23363_/Y sky130_fd_sc_hd__inv_2
X_20575_ _20575_/A vssd1 vssd1 vccd1 vccd1 _20575_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25102_ _27081_/Q _27113_/Q _25102_/S vssd1 vssd1 vccd1 vccd1 _25102_/X sky130_fd_sc_hd__mux2_1
X_22314_ _22314_/A vssd1 vssd1 vccd1 vccd1 _22314_/X sky130_fd_sc_hd__clkbuf_1
X_26082_ _19600_/X _26082_/D vssd1 vssd1 vccd1 vccd1 _26082_/Q sky130_fd_sc_hd__dfxtp_1
X_23294_ _27750_/Q input62/X vssd1 vssd1 vccd1 vccd1 _23300_/A sky130_fd_sc_hd__xor2_1
XFILLER_152_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25033_ _27969_/A _25031_/X _25067_/S vssd1 vssd1 vccd1 vccd1 _25034_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22245_ _22261_/A vssd1 vssd1 vccd1 vccd1 _22245_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22176_ _22176_/A vssd1 vssd1 vccd1 vccd1 _22176_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21127_ _21127_/A vssd1 vssd1 vccd1 vccd1 _21127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26984_ _22750_/X _26984_/D vssd1 vssd1 vccd1 vccd1 _26984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25935_ _25935_/CLK _25935_/D vssd1 vssd1 vccd1 vccd1 _25935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21058_ _21125_/A vssd1 vssd1 vccd1 vccd1 _21058_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20009_ _20076_/A vssd1 vssd1 vccd1 vccd1 _20009_/X sky130_fd_sc_hd__clkbuf_1
X_25866_ _27153_/CLK _25866_/D vssd1 vssd1 vccd1 vccd1 _25866_/Q sky130_fd_sc_hd__dfxtp_1
X_13880_ _13919_/A vssd1 vssd1 vccd1 vccd1 _13880_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27605_ _27606_/CLK _27605_/D vssd1 vssd1 vccd1 vccd1 _27605_/Q sky130_fd_sc_hd__dfxtp_1
X_24817_ _24914_/A vssd1 vssd1 vccd1 vccd1 _24817_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25797_ _17511_/X _27853_/Q _25801_/S vssd1 vssd1 vccd1 vccd1 _25798_/A sky130_fd_sc_hd__mux2_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _15550_/A vssd1 vssd1 vccd1 vccd1 _26202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27536_ _27536_/CLK _27536_/D vssd1 vssd1 vccd1 vccd1 _27536_/Q sky130_fd_sc_hd__dfxtp_2
X_24748_ _24748_/A vssd1 vssd1 vccd1 vccd1 _24940_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _15758_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _14501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27467_ _27467_/CLK _27467_/D vssd1 vssd1 vccd1 vccd1 _27467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15549_/S vssd1 vssd1 vccd1 vccd1 _15490_/S sky130_fd_sc_hd__clkbuf_2
X_24679_ _27173_/Q _24685_/B vssd1 vssd1 vccd1 vccd1 _24679_/X sky130_fd_sc_hd__or2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17220_/A vssd1 vssd1 vccd1 vccd1 _17220_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14432_ _26646_/Q _14421_/X _14416_/X _14431_/Y vssd1 vssd1 vccd1 vccd1 _26646_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26418_ _20767_/X _26418_/D vssd1 vssd1 vccd1 vccd1 _26418_/Q sky130_fd_sc_hd__dfxtp_1
X_27398_ _27398_/CLK _27398_/D vssd1 vssd1 vccd1 vccd1 _27398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17151_ _17149_/X _17150_/X _17174_/S vssd1 vssd1 vccd1 vccd1 _17151_/X sky130_fd_sc_hd__mux2_1
X_14363_ _14363_/A _14363_/B vssd1 vssd1 vccd1 vccd1 _14363_/Y sky130_fd_sc_hd__nor2_1
X_26349_ _20529_/X _26349_/D vssd1 vssd1 vccd1 vccd1 _26349_/Q sky130_fd_sc_hd__dfxtp_1
Xinput16 la1_data_in[16] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_4
XFILLER_168_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 la1_data_in[26] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_4
XFILLER_156_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16102_ _25910_/Q vssd1 vssd1 vccd1 vccd1 _16369_/A sky130_fd_sc_hd__inv_2
Xinput38 la1_data_in[7] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_4
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ _13314_/A vssd1 vssd1 vccd1 vccd1 _27004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput49 la1_oenb[17] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_6
X_17082_ _27832_/Q _27136_/Q _25881_/Q _25849_/Q _17081_/X _17069_/X vssd1 vssd1 vccd1
+ vccd1 _17082_/X sky130_fd_sc_hd__mux4_1
X_14294_ _14383_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14294_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ _16033_/A _16287_/A _16298_/C vssd1 vssd1 vccd1 vccd1 _16033_/X sky130_fd_sc_hd__or3_1
XFILLER_109_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _13672_/B _13425_/A _13672_/A vssd1 vssd1 vccd1 vccd1 _15407_/A sky130_fd_sc_hd__or3b_4
X_28019_ _28019_/A _15984_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
XFILLER_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _27281_/Q _13176_/B vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__and2_1
XFILLER_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17984_ _26271_/Q _26239_/Q _26207_/Q _26175_/Q _17873_/X _17937_/X vssd1 vssd1 vccd1
+ vccd1 _17984_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19723_ _19723_/A vssd1 vssd1 vccd1 vccd1 _19723_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16935_ _27597_/Q _24210_/A _27487_/Q _18443_/A _16934_/X vssd1 vssd1 vccd1 vccd1
+ _16935_/X sky130_fd_sc_hd__o221a_1
XFILLER_78_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19654_ _19637_/X _19638_/X _19639_/X _19640_/X _19644_/X _19647_/X vssd1 vssd1 vccd1
+ vccd1 _19655_/A sky130_fd_sc_hd__mux4_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16866_ _16866_/A _16337_/X vssd1 vssd1 vccd1 vccd1 _16867_/A sky130_fd_sc_hd__or2b_1
XFILLER_19_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18605_ _18605_/A vssd1 vssd1 vccd1 vccd1 _25564_/A sky130_fd_sc_hd__clkbuf_2
X_15817_ _15817_/A vssd1 vssd1 vccd1 vccd1 _26091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19585_ _19570_/X _19572_/X _19574_/X _19576_/X _19577_/X _19578_/X vssd1 vssd1 vccd1
+ vccd1 _19586_/A sky130_fd_sc_hd__mux4_1
X_16797_ _16797_/A _16798_/B vssd1 vssd1 vccd1 vccd1 _16797_/X sky130_fd_sc_hd__or2_1
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18536_ _18009_/X _18533_/X _18535_/X _18014_/X vssd1 vssd1 vccd1 vccd1 _18536_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _15761_/A vssd1 vssd1 vccd1 vccd1 _15758_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _18467_/A vssd1 vssd1 vccd1 vccd1 _25969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_290 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ _15679_/A vssd1 vssd1 vccd1 vccd1 _26145_/D sky130_fd_sc_hd__clkbuf_1
X_17418_ _17418_/A _17418_/B _17418_/C vssd1 vssd1 vccd1 vccd1 _17419_/C sky130_fd_sc_hd__or3_1
XFILLER_21_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18398_ _18398_/A _18398_/B _18398_/C vssd1 vssd1 vccd1 vccd1 _18399_/A sky130_fd_sc_hd__and3_1
XFILLER_140_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17349_ _27854_/Q _27158_/Q _25903_/Q _25871_/Q _17325_/X _17313_/X vssd1 vssd1 vccd1
+ vccd1 _17349_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20360_ _20426_/A vssd1 vssd1 vccd1 vccd1 _20360_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27958__444 vssd1 vssd1 vccd1 vccd1 _27958__444/HI _27958_/A sky130_fd_sc_hd__conb_1
XFILLER_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19019_ _19321_/A vssd1 vssd1 vccd1 vccd1 _19019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20291_ _20323_/A vssd1 vssd1 vccd1 vccd1 _20291_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22030_ _22030_/A vssd1 vssd1 vccd1 vccd1 _22030_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23981_ _27089_/Q _23954_/X _23955_/X _27121_/Q _23956_/X vssd1 vssd1 vccd1 vccd1
+ _23981_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25720_ _25720_/A vssd1 vssd1 vccd1 vccd1 _25720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22932_ _22932_/A vssd1 vssd1 vccd1 vccd1 _22932_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25651_ _25635_/X _25636_/X _25637_/X _25638_/X _25640_/X _25642_/X vssd1 vssd1 vccd1
+ vccd1 _25652_/A sky130_fd_sc_hd__mux4_1
XFILLER_3_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22863_ _22853_/X _22854_/X _22855_/X _22856_/X _22857_/X _22858_/X vssd1 vssd1 vccd1
+ vccd1 _22864_/A sky130_fd_sc_hd__mux4_1
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24602_ _24602_/A vssd1 vssd1 vccd1 vccd1 _27560_/D sky130_fd_sc_hd__clkbuf_1
X_21814_ _21814_/A vssd1 vssd1 vccd1 vccd1 _21814_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25582_ _25582_/A vssd1 vssd1 vccd1 vccd1 _25582_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22794_ _22794_/A vssd1 vssd1 vccd1 vccd1 _22794_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27321_ _27331_/CLK _27321_/D vssd1 vssd1 vccd1 vccd1 _27321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24533_ _24533_/A vssd1 vssd1 vccd1 vccd1 _27532_/D sky130_fd_sc_hd__clkbuf_1
X_21745_ _22089_/A vssd1 vssd1 vccd1 vccd1 _21814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27252_ _27782_/CLK _27252_/D vssd1 vssd1 vccd1 vccd1 _27252_/Q sky130_fd_sc_hd__dfxtp_1
X_24464_ _24464_/A vssd1 vssd1 vccd1 vccd1 _27508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21676_ _21740_/A vssd1 vssd1 vccd1 vccd1 _21676_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_185_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26203_ _20025_/X _26203_/D vssd1 vssd1 vccd1 vccd1 _26203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23415_ _23429_/A vssd1 vssd1 vccd1 vccd1 _23415_/X sky130_fd_sc_hd__clkbuf_2
X_20627_ _20627_/A vssd1 vssd1 vccd1 vccd1 _20627_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27183_ _27601_/CLK _27183_/D vssd1 vssd1 vccd1 vccd1 _27183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24395_ _24395_/A vssd1 vssd1 vccd1 vccd1 _27477_/D sky130_fd_sc_hd__clkbuf_1
X_26134_ _19779_/X _26134_/D vssd1 vssd1 vccd1 vccd1 _26134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23346_ _27778_/Q _27258_/Q vssd1 vssd1 vccd1 vccd1 _23346_/Y sky130_fd_sc_hd__xnor2_1
X_20558_ _20550_/X _20551_/X _20552_/X _20553_/X _20554_/X _20555_/X vssd1 vssd1 vccd1
+ vccd1 _20559_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26065_ _26065_/CLK _26065_/D vssd1 vssd1 vccd1 vccd1 _26065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23277_ _27745_/Q vssd1 vssd1 vccd1 vccd1 _23277_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20489_ _20489_/A vssd1 vssd1 vccd1 vccd1 _20489_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13030_ _13530_/A vssd1 vssd1 vccd1 vccd1 _13030_/X sky130_fd_sc_hd__clkbuf_4
X_25016_ _27967_/A _25015_/X _25024_/S vssd1 vssd1 vccd1 vccd1 _25017_/A sky130_fd_sc_hd__mux2_1
X_22228_ _22228_/A vssd1 vssd1 vccd1 vccd1 _22228_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22159_ _22175_/A vssd1 vssd1 vccd1 vccd1 _22159_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1087 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14981_ _15718_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14981_/Y sky130_fd_sc_hd__nor2_1
X_26967_ _22692_/X _26967_/D vssd1 vssd1 vccd1 vccd1 _26967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16720_ _16722_/A _16786_/B vssd1 vssd1 vccd1 vccd1 _16721_/A sky130_fd_sc_hd__nand2_1
X_13932_ _14172_/A vssd1 vssd1 vccd1 vccd1 _14005_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25918_ _25984_/CLK _25918_/D vssd1 vssd1 vccd1 vccd1 _25918_/Q sky130_fd_sc_hd__dfxtp_1
X_26898_ _22448_/X _26898_/D vssd1 vssd1 vccd1 vccd1 _26898_/Q sky130_fd_sc_hd__dfxtp_1
X_13863_ _15773_/A vssd1 vssd1 vccd1 vccd1 _14172_/A sky130_fd_sc_hd__clkbuf_2
X_16651_ _16651_/A vssd1 vssd1 vccd1 vccd1 _16652_/A sky130_fd_sc_hd__inv_2
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25849_ _25984_/CLK _25849_/D vssd1 vssd1 vccd1 vccd1 _25849_/Q sky130_fd_sc_hd__dfxtp_1
X_15602_ _26179_/Q _16235_/A _15606_/S vssd1 vssd1 vccd1 vccd1 _15603_/A sky130_fd_sc_hd__mux2_1
X_19370_ _26832_/Q _26800_/Q _26768_/Q _26736_/Q _18913_/X _18930_/X vssd1 vssd1 vccd1
+ vccd1 _19370_/X sky130_fd_sc_hd__mux4_2
X_13794_ _13833_/A vssd1 vssd1 vccd1 vccd1 _13794_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16582_ _16576_/A _16561_/A _16561_/B vssd1 vssd1 vccd1 vccd1 _16583_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18321_ _26157_/Q _26093_/Q _27021_/Q _26989_/Q _18298_/X _18228_/X vssd1 vssd1 vccd1
+ vccd1 _18323_/A sky130_fd_sc_hd__mux4_1
X_15533_ _15533_/A vssd1 vssd1 vccd1 vccd1 _26210_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27519_ _27574_/CLK _27519_/D vssd1 vssd1 vccd1 vccd1 _27519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18252_ _18198_/X _18248_/X _18251_/X _18203_/X vssd1 vssd1 vccd1 vccd1 _18252_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15464_ _15464_/A vssd1 vssd1 vccd1 vccd1 _15473_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17203_ _17325_/A vssd1 vssd1 vccd1 vccd1 _17203_/X sky130_fd_sc_hd__buf_2
X_14415_ _14436_/A vssd1 vssd1 vccd1 vccd1 _14532_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15395_ _14795_/X _26271_/Q _15401_/S vssd1 vssd1 vccd1 vccd1 _15396_/A sky130_fd_sc_hd__mux2_1
X_18183_ _26151_/Q _26087_/Q _27015_/Q _26983_/Q _18182_/X _18112_/X vssd1 vssd1 vccd1
+ vccd1 _18184_/A sky130_fd_sc_hd__mux4_1
XFILLER_129_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14346_ _14346_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _14346_/Y sky130_fd_sc_hd__nor2_1
X_17134_ _25821_/Q _26020_/Q _17158_/S vssd1 vssd1 vccd1 vccd1 _17134_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _17386_/S vssd1 vssd1 vccd1 vccd1 _17113_/S sky130_fd_sc_hd__clkbuf_2
X_14277_ _26701_/Q _14270_/X _14271_/X _14276_/Y vssd1 vssd1 vccd1 vccd1 _26701_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_195_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16016_ _27482_/Q _27269_/Q vssd1 vssd1 vccd1 vccd1 _16016_/X sky130_fd_sc_hd__or2_1
X_13228_ _14804_/A vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__buf_2
XFILLER_170_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13159_ _27284_/Q _13176_/B vssd1 vssd1 vccd1 vccd1 _13159_/X sky130_fd_sc_hd__and2_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _18405_/A vssd1 vssd1 vccd1 vccd1 _18075_/S sky130_fd_sc_hd__clkbuf_2
Xrepeater403 _27365_/CLK vssd1 vssd1 vccd1 vccd1 _27357_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater414 _27334_/CLK vssd1 vssd1 vccd1 vccd1 _27311_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater425 _26056_/CLK vssd1 vssd1 vccd1 vccd1 _26057_/CLK sky130_fd_sc_hd__clkbuf_1
X_19706_ _19694_/X _19695_/X _19696_/X _19697_/X _19698_/X _19699_/X vssd1 vssd1 vccd1
+ vccd1 _19707_/A sky130_fd_sc_hd__mux4_1
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16918_ _16833_/A _16916_/Y _16917_/X vssd1 vssd1 vccd1 vccd1 _16918_/X sky130_fd_sc_hd__o21a_1
X_17898_ _17898_/A vssd1 vssd1 vccd1 vccd1 _18462_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19637_ _19637_/A vssd1 vssd1 vccd1 vccd1 _19637_/X sky130_fd_sc_hd__clkbuf_1
X_16849_ _16200_/B _16759_/B _16848_/X vssd1 vssd1 vccd1 vccd1 _16849_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19568_ _19568_/A vssd1 vssd1 vccd1 vccd1 _26073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18519_ _17897_/X _18514_/X _18516_/X _18518_/X _18352_/S vssd1 vssd1 vccd1 vccd1
+ _18528_/B sky130_fd_sc_hd__a221o_1
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19499_ _19497_/X _19498_/X _19499_/S vssd1 vssd1 vccd1 vccd1 _19499_/X sky130_fd_sc_hd__mux2_1
X_21530_ _21562_/A vssd1 vssd1 vccd1 vccd1 _21530_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21461_ _21477_/A vssd1 vssd1 vccd1 vccd1 _21461_/X sky130_fd_sc_hd__clkbuf_1
X_23200_ _17447_/X _27137_/Q _23204_/S vssd1 vssd1 vccd1 vccd1 _23201_/A sky130_fd_sc_hd__mux2_1
X_20412_ _20412_/A vssd1 vssd1 vccd1 vccd1 _20412_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24180_ _27466_/Q _24184_/B vssd1 vssd1 vccd1 vccd1 _24181_/A sky130_fd_sc_hd__and2_1
X_21392_ _21392_/A vssd1 vssd1 vccd1 vccd1 _21392_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23131_ _23131_/A vssd1 vssd1 vccd1 vccd1 _27106_/D sky130_fd_sc_hd__clkbuf_1
X_20343_ _20343_/A vssd1 vssd1 vccd1 vccd1 _20343_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_179_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23062_ _27076_/Q _17708_/X _23070_/S vssd1 vssd1 vccd1 vccd1 _23063_/A sky130_fd_sc_hd__mux2_1
X_20274_ _20322_/A vssd1 vssd1 vccd1 vccd1 _20274_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22013_ _21997_/X _21998_/X _21999_/X _22000_/X _22002_/X _22004_/X vssd1 vssd1 vccd1
+ vccd1 _22014_/A sky130_fd_sc_hd__mux4_1
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26821_ _22186_/X _26821_/D vssd1 vssd1 vccd1 vccd1 _26821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26752_ _21944_/X _26752_/D vssd1 vssd1 vccd1 vccd1 _26752_/Q sky130_fd_sc_hd__dfxtp_1
X_23964_ _23962_/X _23963_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23964_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_6 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25703_ _25689_/X _25690_/X _25691_/X _25692_/X _25693_/X _25694_/X vssd1 vssd1 vccd1
+ vccd1 _25704_/A sky130_fd_sc_hd__mux4_1
XFILLER_56_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22915_ _22907_/X _22908_/X _22909_/X _22910_/X _22911_/X _22912_/X vssd1 vssd1 vccd1
+ vccd1 _22916_/A sky130_fd_sc_hd__mux4_1
X_26683_ _21702_/X _26683_/D vssd1 vssd1 vccd1 vccd1 _26683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23895_ _23849_/X _23893_/X _23894_/X _23864_/X vssd1 vssd1 vccd1 vccd1 _27285_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22846_ _22846_/A vssd1 vssd1 vccd1 vccd1 _22846_/X sky130_fd_sc_hd__clkbuf_1
X_25634_ _25634_/A vssd1 vssd1 vccd1 vccd1 _25634_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25565_ _25547_/X _25552_/X _25553_/X _24928_/B _25554_/X vssd1 vssd1 vccd1 vccd1
+ _25565_/X sky130_fd_sc_hd__o311a_1
XFILLER_169_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22777_ _22767_/X _22768_/X _22769_/X _22770_/X _22771_/X _22772_/X vssd1 vssd1 vccd1
+ vccd1 _22778_/A sky130_fd_sc_hd__mux4_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24516_ _24516_/A vssd1 vssd1 vccd1 vccd1 _27527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27304_ _27377_/CLK _27304_/D vssd1 vssd1 vccd1 vccd1 _27304_/Q sky130_fd_sc_hd__dfxtp_1
X_21728_ _21728_/A vssd1 vssd1 vccd1 vccd1 _21728_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25496_ _25470_/X _25192_/B _25495_/X _25483_/X vssd1 vssd1 vccd1 vccd1 _25496_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24447_ _24480_/A vssd1 vssd1 vccd1 vccd1 _24456_/B sky130_fd_sc_hd__clkbuf_1
X_27235_ _27236_/CLK _27235_/D vssd1 vssd1 vccd1 vccd1 _27235_/Q sky130_fd_sc_hd__dfxtp_1
X_21659_ _21647_/X _21648_/X _21649_/X _21650_/X _21652_/X _21654_/X vssd1 vssd1 vccd1
+ vccd1 _21660_/A sky130_fd_sc_hd__mux4_1
X_14200_ _14376_/A _14200_/B vssd1 vssd1 vccd1 vccd1 _14200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15180_ _26366_/Q _13408_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15181_/A sky130_fd_sc_hd__mux2_1
X_27166_ _27578_/CLK _27166_/D vssd1 vssd1 vccd1 vccd1 _27166_/Q sky130_fd_sc_hd__dfxtp_1
X_24378_ _27571_/Q _24380_/B vssd1 vssd1 vccd1 vccd1 _24379_/A sky130_fd_sc_hd__and2_1
XFILLER_138_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14131_ _14396_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14131_/Y sky130_fd_sc_hd__nor2_1
X_26117_ _19721_/X _26117_/D vssd1 vssd1 vccd1 vccd1 _26117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23329_ input48/X input49/X input50/X input51/X vssd1 vssd1 vccd1 vccd1 _23331_/C
+ sky130_fd_sc_hd__or4_1
X_27097_ _27109_/CLK _27097_/D vssd1 vssd1 vccd1 vccd1 _27097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14062_ _15190_/A _14149_/B vssd1 vssd1 vccd1 vccd1 _14079_/A sky130_fd_sc_hd__or2_1
XFILLER_125_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26048_ _26048_/CLK _26048_/D vssd1 vssd1 vccd1 vccd1 _26048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ _27793_/Q _25733_/B vssd1 vssd1 vccd1 vccd1 _13014_/A sky130_fd_sc_hd__and2_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18870_ _19338_/A vssd1 vssd1 vccd1 vccd1 _18870_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17821_ _18182_/A vssd1 vssd1 vccd1 vccd1 _17821_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27999_ _27999_/A _15881_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
XFILLER_43_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17752_ _17752_/A vssd1 vssd1 vccd1 vccd1 _25935_/D sky130_fd_sc_hd__clkbuf_1
X_14964_ _15701_/A _14966_/B vssd1 vssd1 vccd1 vccd1 _14964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16703_ _16703_/A _16703_/B vssd1 vssd1 vccd1 vccd1 _16703_/X sky130_fd_sc_hd__xor2_1
X_13915_ _13915_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _13915_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17683_ _27410_/Q vssd1 vssd1 vccd1 vccd1 _17683_/X sky130_fd_sc_hd__clkbuf_2
X_14895_ _14895_/A vssd1 vssd1 vccd1 vccd1 _26486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19422_ _26418_/Q _26386_/Q _26354_/Q _26322_/Q _19331_/X _19399_/X vssd1 vssd1 vccd1
+ vccd1 _19422_/X sky130_fd_sc_hd__mux4_1
X_16634_ _16621_/X _16807_/B _16807_/A vssd1 vssd1 vccd1 vccd1 _16634_/X sky130_fd_sc_hd__o21ba_1
X_13846_ _26843_/Q _13844_/X _13770_/B _13845_/Y vssd1 vssd1 vccd1 vccd1 _26843_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19353_ _26287_/Q _26255_/Q _26223_/Q _26191_/Q _19283_/X _19352_/X vssd1 vssd1 vccd1
+ vccd1 _19353_/X sky130_fd_sc_hd__mux4_1
X_13777_ _26869_/Q _13761_/X _13764_/X _13776_/Y vssd1 vssd1 vccd1 vccd1 _26869_/D
+ sky130_fd_sc_hd__a31o_1
X_16565_ _16565_/A vssd1 vssd1 vccd1 vccd1 _16798_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18304_ _26540_/Q _26508_/Q _26476_/Q _27052_/Q _18233_/X _18259_/X vssd1 vssd1 vccd1
+ vccd1 _18304_/X sky130_fd_sc_hd__mux4_1
X_15516_ _15516_/A vssd1 vssd1 vccd1 vccd1 _26218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19284_ _26284_/Q _26252_/Q _26220_/Q _26188_/Q _19283_/X _19192_/X vssd1 vssd1 vccd1
+ vccd1 _19284_/X sky130_fd_sc_hd__mux4_1
X_16496_ _27392_/Q _16094_/X _16098_/X _25960_/Q _16495_/Y vssd1 vssd1 vccd1 vccd1
+ _16499_/A sky130_fd_sc_hd__a221oi_4
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18235_ _26409_/Q _26377_/Q _26345_/Q _26313_/Q _18189_/X _18214_/X vssd1 vssd1 vccd1
+ vccd1 _18235_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15447_ _26248_/Q _13376_/X _15451_/S vssd1 vssd1 vccd1 vccd1 _15448_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18166_ _26406_/Q _26374_/Q _26342_/Q _26310_/Q _18048_/X _18073_/X vssd1 vssd1 vccd1
+ vccd1 _18166_/X sky130_fd_sc_hd__mux4_1
XFILLER_172_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15378_ _15378_/A vssd1 vssd1 vccd1 vccd1 _26279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _27835_/Q _27139_/Q _25884_/Q _25852_/Q _17081_/X _17069_/X vssd1 vssd1 vccd1
+ vccd1 _17117_/X sky130_fd_sc_hd__mux4_1
X_14329_ _14412_/B vssd1 vssd1 vccd1 vccd1 _14329_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18097_ _18146_/A _18097_/B _18097_/C vssd1 vssd1 vccd1 vccd1 _18098_/A sky130_fd_sc_hd__and3_1
XFILLER_172_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17048_ _17046_/X _17047_/X _17048_/S vssd1 vssd1 vccd1 vccd1 _17048_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_509 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater200 _25923_/CLK vssd1 vssd1 vccd1 vccd1 _27141_/CLK sky130_fd_sc_hd__clkbuf_1
X_18999_ _26944_/Q _26912_/Q _26880_/Q _26848_/Q _18875_/X _18972_/X vssd1 vssd1 vccd1
+ vccd1 _18999_/X sky130_fd_sc_hd__mux4_2
Xrepeater211 _27076_/CLK vssd1 vssd1 vccd1 vccd1 _25913_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater222 _27406_/CLK vssd1 vssd1 vccd1 vccd1 _27404_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater233 _27735_/CLK vssd1 vssd1 vccd1 vccd1 _27750_/CLK sky130_fd_sc_hd__clkbuf_2
Xrepeater244 _27749_/CLK vssd1 vssd1 vccd1 vccd1 _27623_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater255 _27614_/CLK vssd1 vssd1 vccd1 vccd1 _27617_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater266 _27593_/CLK vssd1 vssd1 vccd1 vccd1 _27172_/CLK sky130_fd_sc_hd__clkbuf_1
X_20961_ _20953_/X _20954_/X _20955_/X _20956_/X _20958_/X _20960_/X vssd1 vssd1 vccd1
+ vccd1 _20962_/A sky130_fd_sc_hd__mux4_1
Xrepeater277 _27610_/CLK vssd1 vssd1 vccd1 vccd1 _27539_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater288 _27478_/CLK vssd1 vssd1 vccd1 vccd1 _27477_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater299 _27649_/CLK vssd1 vssd1 vccd1 vccd1 _27236_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22700_ _22700_/A vssd1 vssd1 vccd1 vccd1 _22700_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23680_ _23680_/A vssd1 vssd1 vccd1 vccd1 _27245_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20892_ _20956_/A vssd1 vssd1 vccd1 vccd1 _20892_/X sky130_fd_sc_hd__clkbuf_1
X_22631_ _22889_/A vssd1 vssd1 vccd1 vccd1 _22698_/A sky130_fd_sc_hd__buf_2
XFILLER_81_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25350_ _25350_/A _25350_/B vssd1 vssd1 vccd1 vccd1 _25351_/B sky130_fd_sc_hd__xnor2_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22562_ _22610_/A vssd1 vssd1 vccd1 vccd1 _22562_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24301_ _24301_/A _24302_/B vssd1 vssd1 vccd1 vccd1 _27431_/D sky130_fd_sc_hd__nor2_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21513_ _21561_/A vssd1 vssd1 vccd1 vccd1 _21513_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25281_ _25354_/A _27507_/Q _25273_/A vssd1 vssd1 vccd1 vccd1 _25282_/B sky130_fd_sc_hd__a21o_1
X_22493_ _22487_/X _22488_/X _22489_/X _22490_/X _22491_/X _22492_/X vssd1 vssd1 vccd1
+ vccd1 _22494_/A sky130_fd_sc_hd__mux4_1
XFILLER_186_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27020_ _22878_/X _27020_/D vssd1 vssd1 vccd1 vccd1 _27020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24232_ _24232_/A _24235_/B vssd1 vssd1 vccd1 vccd1 _27387_/D sky130_fd_sc_hd__nor2_1
X_21444_ _21476_/A vssd1 vssd1 vccd1 vccd1 _21444_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24163_ _24163_/A vssd1 vssd1 vccd1 vccd1 _27353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21375_ _21391_/A vssd1 vssd1 vccd1 vccd1 _21375_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23114_ _23114_/A vssd1 vssd1 vccd1 vccd1 _27098_/D sky130_fd_sc_hd__clkbuf_1
X_20326_ _20318_/X _20319_/X _20320_/X _20321_/X _20322_/X _20323_/X vssd1 vssd1 vccd1
+ vccd1 _20327_/A sky130_fd_sc_hd__mux4_1
X_24094_ _24094_/A vssd1 vssd1 vccd1 vccd1 _27322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27922_ _27922_/A _15965_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
X_23045_ _23045_/A vssd1 vssd1 vccd1 vccd1 _27068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20257_ _20257_/A vssd1 vssd1 vccd1 vccd1 _20257_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_658 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27853_ _27855_/CLK _27853_/D vssd1 vssd1 vccd1 vccd1 _27853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20188_ _20236_/A vssd1 vssd1 vccd1 vccd1 _20188_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26804_ _22124_/X _26804_/D vssd1 vssd1 vccd1 vccd1 _26804_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27784_ _27784_/CLK _27784_/D vssd1 vssd1 vccd1 vccd1 _27784_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24996_ _27232_/Q vssd1 vssd1 vccd1 vccd1 _25103_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26735_ _21886_/X _26735_/D vssd1 vssd1 vccd1 vccd1 _26735_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23947_ _25932_/Q _25998_/Q _25831_/Q _26030_/Q _23946_/X _23929_/X vssd1 vssd1 vccd1
+ vccd1 _23947_/X sky130_fd_sc_hd__mux4_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _13740_/A vssd1 vssd1 vccd1 vccd1 _13711_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _15754_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26666_ _21640_/X _26666_/D vssd1 vssd1 vccd1 vccd1 _26666_/Q sky130_fd_sc_hd__dfxtp_1
X_23878_ _23876_/X _23877_/X _23893_/S vssd1 vssd1 vccd1 vccd1 _23878_/X sky130_fd_sc_hd__mux2_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ _26922_/Q _13626_/X _13629_/X _13630_/Y vssd1 vssd1 vccd1 vccd1 _26922_/D
+ sky130_fd_sc_hd__a31o_1
X_25617_ _25617_/A _25618_/B vssd1 vssd1 vccd1 vccd1 _27787_/D sky130_fd_sc_hd__nor2_1
X_22829_ _22821_/X _22822_/X _22823_/X _22824_/X _22825_/X _22826_/X vssd1 vssd1 vccd1
+ vccd1 _22830_/A sky130_fd_sc_hd__mux4_1
X_26597_ _21402_/X _26597_/D vssd1 vssd1 vccd1 vccd1 _26597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13562_ _26943_/Q _13558_/X _13553_/X _13561_/Y vssd1 vssd1 vccd1 vccd1 _26943_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16350_ _16337_/X _16867_/B _16866_/A vssd1 vssd1 vccd1 vccd1 _16858_/B sky130_fd_sc_hd__a21o_1
X_25548_ _25547_/X _25522_/X _25523_/X _24913_/B _25524_/X vssd1 vssd1 vccd1 vccd1
+ _25548_/X sky130_fd_sc_hd__o311a_1
XFILLER_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15301_ _15301_/A vssd1 vssd1 vccd1 vccd1 _26313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16281_ _16633_/A _16281_/B vssd1 vssd1 vccd1 vccd1 _16292_/C sky130_fd_sc_hd__or2_1
X_13493_ _14464_/A vssd1 vssd1 vccd1 vccd1 _13891_/A sky130_fd_sc_hd__clkbuf_2
X_25479_ _25539_/A vssd1 vssd1 vccd1 vccd1 _25479_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18020_ _18020_/A vssd1 vssd1 vccd1 vccd1 _18020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27218_ _27422_/CLK _27218_/D vssd1 vssd1 vccd1 vccd1 _27218_/Q sky130_fd_sc_hd__dfxtp_1
X_15232_ _14769_/X _26343_/Q _15234_/S vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _15163_/A vssd1 vssd1 vccd1 vccd1 _26374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27149_ _27149_/CLK _27149_/D vssd1 vssd1 vccd1 vccd1 _27149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14114_ _14127_/A vssd1 vssd1 vccd1 vccd1 _14125_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ _15094_/A vssd1 vssd1 vccd1 vccd1 _26405_/D sky130_fd_sc_hd__clkbuf_1
X_19971_ _19971_/A vssd1 vssd1 vccd1 vccd1 _19971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14045_ _26783_/Q _14042_/X _14038_/X _14044_/Y vssd1 vssd1 vccd1 vccd1 _26783_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_140_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18922_ _18922_/A vssd1 vssd1 vccd1 vccd1 _18922_/X sky130_fd_sc_hd__buf_4
XFILLER_140_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18853_ _18850_/X _18852_/X _19560_/A vssd1 vssd1 vccd1 vccd1 _18853_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_28015__481 vssd1 vssd1 vccd1 vccd1 _28015__481/HI _28015_/A sky130_fd_sc_hd__conb_1
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17804_ _18000_/A vssd1 vssd1 vccd1 vccd1 _18012_/A sky130_fd_sc_hd__clkbuf_2
X_18784_ _27601_/Q vssd1 vssd1 vccd1 vccd1 _18932_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15996_ _16593_/A vssd1 vssd1 vccd1 vccd1 _16623_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17735_ _25930_/Q _17734_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17736_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14947_ _14798_/X _26462_/Q _14951_/S vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17666_ _17666_/A vssd1 vssd1 vccd1 vccd1 _25903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14878_ _14878_/A vssd1 vssd1 vccd1 vccd1 _26493_/D sky130_fd_sc_hd__clkbuf_1
X_19405_ _19471_/A _19405_/B _19405_/C vssd1 vssd1 vccd1 vccd1 _19406_/A sky130_fd_sc_hd__and3_1
X_16617_ _16614_/Y _16885_/B _16616_/X vssd1 vssd1 vccd1 vccd1 _16618_/B sky130_fd_sc_hd__o21bai_1
X_13829_ _26850_/Q _13819_/X _13820_/X _13828_/Y vssd1 vssd1 vccd1 vccd1 _26850_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17597_ _17520_/X _25873_/Q _17599_/S vssd1 vssd1 vccd1 vccd1 _17598_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19336_ _19362_/A _19336_/B _19336_/C vssd1 vssd1 vccd1 vccd1 _19337_/A sky130_fd_sc_hd__and3_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16548_ _16535_/A _16535_/B _16547_/X vssd1 vssd1 vccd1 vccd1 _16548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19267_ _19261_/X _19263_/X _19266_/X _19151_/X _19220_/X vssd1 vssd1 vccd1 vccd1
+ _19268_/C sky130_fd_sc_hd__a221o_1
X_16479_ _16479_/A _16479_/B vssd1 vssd1 vccd1 vccd1 _16479_/Y sky130_fd_sc_hd__nand2_1
X_18218_ _18264_/A _18218_/B _18218_/C vssd1 vssd1 vccd1 vccd1 _18219_/A sky130_fd_sc_hd__and3_1
XFILLER_148_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19198_ _19492_/A vssd1 vssd1 vccd1 vccd1 _19334_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18149_ _18844_/A vssd1 vssd1 vccd1 vccd1 _18264_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_117_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21160_ _21160_/A vssd1 vssd1 vccd1 vccd1 _21160_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20111_ _20111_/A vssd1 vssd1 vccd1 vccd1 _20111_/X sky130_fd_sc_hd__clkbuf_1
X_21091_ _21077_/X _21078_/X _21079_/X _21080_/X _21081_/X _21082_/X vssd1 vssd1 vccd1
+ vccd1 _21092_/A sky130_fd_sc_hd__mux4_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20042_ _20028_/X _20029_/X _20030_/X _20031_/X _20032_/X _20033_/X vssd1 vssd1 vccd1
+ vccd1 _20043_/A sky130_fd_sc_hd__mux4_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24850_ _27646_/Q _24834_/X _24849_/Y _24839_/X vssd1 vssd1 vccd1 vccd1 _27646_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23801_ _27786_/Q vssd1 vssd1 vccd1 vccd1 _23991_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24781_ _27626_/Q _24771_/X _24780_/Y _24773_/X vssd1 vssd1 vccd1 vccd1 _27626_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21993_ _21981_/X _21982_/X _21983_/X _21984_/X _21985_/X _21986_/X vssd1 vssd1 vccd1
+ vccd1 _21994_/A sky130_fd_sc_hd__mux4_1
XFILLER_113_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _22613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23732_ _27372_/Q _24050_/B vssd1 vssd1 vccd1 vccd1 _23733_/A sky130_fd_sc_hd__and2_1
XFILLER_82_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26520_ _21134_/X _26520_/D vssd1 vssd1 vccd1 vccd1 _26520_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_119 _22546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20944_ _20944_/A vssd1 vssd1 vccd1 vccd1 _20944_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26451_ _20898_/X _26451_/D vssd1 vssd1 vccd1 vccd1 _26451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23663_ _23720_/S vssd1 vssd1 vccd1 vccd1 _23672_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_198_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20875_ _20864_/X _20865_/X _20866_/X _20867_/X _20870_/X _20874_/X vssd1 vssd1 vccd1
+ vccd1 _20876_/A sky130_fd_sc_hd__mux4_1
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22614_ _22959_/A vssd1 vssd1 vccd1 vccd1 _22685_/A sky130_fd_sc_hd__buf_2
X_25402_ _27740_/Q input51/X _25402_/S vssd1 vssd1 vccd1 vccd1 _25403_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26382_ _20647_/X _26382_/D vssd1 vssd1 vccd1 vccd1 _26382_/Q sky130_fd_sc_hd__dfxtp_1
X_23594_ _27777_/Q vssd1 vssd1 vccd1 vccd1 _25580_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_201_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_821 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25333_ _25319_/C _25329_/X _25330_/Y _25331_/Y _25332_/X vssd1 vssd1 vccd1 vccd1
+ _25339_/B sky130_fd_sc_hd__a311o_1
X_22545_ _22611_/A vssd1 vssd1 vccd1 vccd1 _22545_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25264_ _25309_/A vssd1 vssd1 vccd1 vccd1 _25306_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22476_ _22508_/A vssd1 vssd1 vccd1 vccd1 _22476_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24215_ _24215_/A _24233_/B vssd1 vssd1 vccd1 vccd1 _24216_/A sky130_fd_sc_hd__and2_1
X_27003_ _22818_/X _27003_/D vssd1 vssd1 vccd1 vccd1 _27003_/Q sky130_fd_sc_hd__dfxtp_1
X_21427_ _21475_/A vssd1 vssd1 vccd1 vccd1 _21427_/X sky130_fd_sc_hd__clkbuf_1
X_25195_ _27530_/Q _27498_/Q vssd1 vssd1 vccd1 vccd1 _25197_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24146_ _24146_/A vssd1 vssd1 vccd1 vccd1 _27345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21358_ _21390_/A vssd1 vssd1 vccd1 vccd1 _21358_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20309_ _20309_/A vssd1 vssd1 vccd1 vccd1 _20309_/X sky130_fd_sc_hd__clkbuf_1
X_24077_ _24077_/A vssd1 vssd1 vccd1 vccd1 _27314_/D sky130_fd_sc_hd__clkbuf_1
X_21289_ _21289_/A vssd1 vssd1 vccd1 vccd1 _21289_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23028_ _25638_/A vssd1 vssd1 vccd1 vccd1 _23028_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27836_ _27837_/CLK _27836_/D vssd1 vssd1 vccd1 vccd1 _27836_/Q sky130_fd_sc_hd__dfxtp_1
X_15850_ _15850_/A vssd1 vssd1 vccd1 vccd1 _26076_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _14801_/A vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__clkbuf_2
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _15781_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15781_/Y sky130_fd_sc_hd__nor2_1
X_27767_ _27774_/CLK _27767_/D vssd1 vssd1 vccd1 vccd1 _27767_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24979_ _24977_/X _24978_/X _24987_/S vssd1 vssd1 vccd1 vccd1 _24979_/X sky130_fd_sc_hd__mux2_1
X_12993_ _12993_/A vssd1 vssd1 vccd1 vccd1 _27802_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _27438_/Q vssd1 vssd1 vccd1 vccd1 _17520_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26718_ _21822_/X _26718_/D vssd1 vssd1 vccd1 vccd1 _26718_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _14731_/X _26547_/Q _14741_/S vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__mux2_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27698_ _27700_/CLK _27698_/D vssd1 vssd1 vccd1 vccd1 _27698_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17450_/X _25819_/Q _17454_/S vssd1 vssd1 vccd1 vccd1 _17452_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26649_ _21578_/X _26649_/D vssd1 vssd1 vccd1 vccd1 _26649_/Q sky130_fd_sc_hd__dfxtp_1
X_14663_ _26572_/Q _14658_/X _14653_/X _14662_/Y vssd1 vssd1 vccd1 vccd1 _26572_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _16402_/A vssd1 vssd1 vccd1 vccd1 _16557_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13614_ _13884_/A _13621_/B vssd1 vssd1 vccd1 vccd1 _13614_/Y sky130_fd_sc_hd__nor2_1
X_17382_ _25842_/Q _26041_/Q _17382_/S vssd1 vssd1 vccd1 vccd1 _17382_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14594_ _26597_/Q _14589_/X _14592_/X _14593_/Y vssd1 vssd1 vccd1 vccd1 _26597_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19121_ _19113_/X _19115_/X _19120_/X _19022_/X _19023_/X vssd1 vssd1 vccd1 vccd1
+ _19130_/B sky130_fd_sc_hd__a221o_1
X_16333_ _23182_/B _16490_/B vssd1 vssd1 vccd1 vccd1 _16333_/Y sky130_fd_sc_hd__nor2_1
X_13545_ _14503_/A vssd1 vssd1 vccd1 vccd1 _13921_/A sky130_fd_sc_hd__buf_2
XFILLER_41_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19052_ _26274_/Q _26242_/Q _26210_/Q _26178_/Q _19028_/X _18955_/X vssd1 vssd1 vccd1
+ vccd1 _19052_/X sky130_fd_sc_hd__mux4_2
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _13882_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13476_/Y sky130_fd_sc_hd__nor2_1
X_16264_ _27392_/Q _16264_/B vssd1 vssd1 vccd1 vccd1 _16264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_770 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_792 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18003_ _17998_/X _18001_/X _18580_/S vssd1 vssd1 vccd1 vccd1 _18003_/X sky130_fd_sc_hd__mux2_1
X_15215_ _14743_/X _26351_/Q _15223_/S vssd1 vssd1 vccd1 vccd1 _15216_/A sky130_fd_sc_hd__mux2_1
X_16195_ _27379_/Q vssd1 vssd1 vccd1 vccd1 _17410_/A sky130_fd_sc_hd__clkinv_2
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15146_ _15146_/A vssd1 vssd1 vccd1 vccd1 _26382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19954_ _19940_/X _19941_/X _19942_/X _19943_/X _19944_/X _19945_/X vssd1 vssd1 vccd1
+ vccd1 _19955_/A sky130_fd_sc_hd__mux4_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15077_ _14753_/X _26412_/Q _15079_/S vssd1 vssd1 vccd1 vccd1 _15078_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ _14500_/A vssd1 vssd1 vccd1 vccd1 _14390_/A sky130_fd_sc_hd__buf_2
X_18905_ _19296_/S vssd1 vssd1 vccd1 vccd1 _19431_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19885_ _19901_/A vssd1 vssd1 vccd1 vccd1 _19885_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18836_ _19448_/A vssd1 vssd1 vccd1 vccd1 _19290_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18767_ _19338_/A vssd1 vssd1 vccd1 vccd1 _18767_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15979_ _15979_/A vssd1 vssd1 vccd1 vccd1 _15979_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17718_ _27421_/Q vssd1 vssd1 vccd1 vccd1 _17718_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18698_ _26012_/Q _17683_/X _18702_/S vssd1 vssd1 vccd1 vccd1 _18699_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17649_ _17649_/A vssd1 vssd1 vccd1 vccd1 _25895_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20660_ _20652_/X _20653_/X _20654_/X _20655_/X _20656_/X _20657_/X vssd1 vssd1 vccd1
+ vccd1 _20661_/A sky130_fd_sc_hd__mux4_1
XFILLER_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19319_ _19273_/X _19318_/X _19229_/X vssd1 vssd1 vccd1 vccd1 _19319_/X sky130_fd_sc_hd__o21a_1
X_20591_ _20591_/A vssd1 vssd1 vccd1 vccd1 _20591_/X sky130_fd_sc_hd__clkbuf_1
X_22330_ _22330_/A vssd1 vssd1 vccd1 vccd1 _22330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22261_ _22261_/A vssd1 vssd1 vccd1 vccd1 _22261_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24000_ _23996_/X _23998_/X _24033_/S vssd1 vssd1 vccd1 vccd1 _24000_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21212_ _21212_/A vssd1 vssd1 vccd1 vccd1 _21212_/X sky130_fd_sc_hd__clkbuf_1
X_22192_ _22192_/A vssd1 vssd1 vccd1 vccd1 _22192_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21143_ _21143_/A vssd1 vssd1 vccd1 vccd1 _21211_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21074_ _21074_/A vssd1 vssd1 vccd1 vccd1 _21074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25951_ _25953_/CLK _25951_/D vssd1 vssd1 vccd1 vccd1 _25951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24902_ _27770_/Q _24902_/B vssd1 vssd1 vccd1 vccd1 _24903_/B sky130_fd_sc_hd__nor2_1
X_20025_ _20025_/A vssd1 vssd1 vccd1 vccd1 _20025_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25882_ _27833_/CLK _25882_/D vssd1 vssd1 vccd1 vccd1 _25882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27621_ _27621_/CLK _27621_/D vssd1 vssd1 vccd1 vccd1 _27621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24833_ _27643_/Q _24813_/X _24832_/Y _24817_/X vssd1 vssd1 vccd1 vccd1 _27643_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27552_ _27555_/CLK _27552_/D vssd1 vssd1 vccd1 vccd1 _27552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _21976_/A vssd1 vssd1 vccd1 vccd1 _21976_/X sky130_fd_sc_hd__clkbuf_1
X_24764_ _27619_/Q _24758_/X _24763_/Y _24760_/X vssd1 vssd1 vccd1 vccd1 _27619_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26503_ _21074_/X _26503_/D vssd1 vssd1 vccd1 vccd1 _26503_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23715_ _23715_/A vssd1 vssd1 vccd1 vccd1 _27261_/D sky130_fd_sc_hd__clkbuf_1
X_20927_ _20921_/X _20922_/X _20923_/X _20924_/X _20925_/X _20926_/X vssd1 vssd1 vccd1
+ vccd1 _20928_/A sky130_fd_sc_hd__mux4_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24695_ _24392_/A _24687_/X _24694_/X _24690_/X vssd1 vssd1 vccd1 vccd1 _27595_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27483_ _27484_/CLK _27483_/D vssd1 vssd1 vccd1 vccd1 _27483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26434_ _20831_/X _26434_/D vssd1 vssd1 vccd1 vccd1 _26434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20858_ _20848_/X _20849_/X _20850_/X _20851_/X _20852_/X _20853_/X vssd1 vssd1 vccd1
+ vccd1 _20859_/A sky130_fd_sc_hd__mux4_1
X_23646_ _27232_/Q vssd1 vssd1 vccd1 vccd1 _24987_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23577_ _23577_/A _23577_/B vssd1 vssd1 vccd1 vccd1 _23578_/A sky130_fd_sc_hd__and2_1
X_26365_ _20589_/X _26365_/D vssd1 vssd1 vccd1 vccd1 _26365_/Q sky130_fd_sc_hd__dfxtp_1
X_20789_ _22537_/A vssd1 vssd1 vccd1 vccd1 _21143_/A sky130_fd_sc_hd__clkbuf_2
X_13330_ _13330_/A vssd1 vssd1 vccd1 vccd1 _26999_/D sky130_fd_sc_hd__clkbuf_1
X_22528_ _22528_/A vssd1 vssd1 vccd1 vccd1 _22528_/X sky130_fd_sc_hd__clkbuf_1
X_25316_ _27512_/Q _27511_/Q _25332_/A vssd1 vssd1 vccd1 vccd1 _25319_/C sky130_fd_sc_hd__o21ai_1
XFILLER_194_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26296_ _20345_/X _26296_/D vssd1 vssd1 vccd1 vccd1 _26296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _27028_/Q _13086_/X _13269_/S vssd1 vssd1 vccd1 vccd1 _13262_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22459_ _22507_/A vssd1 vssd1 vccd1 vccd1 _22459_/X sky130_fd_sc_hd__clkbuf_2
X_25247_ _27537_/Q _27505_/Q vssd1 vssd1 vccd1 vccd1 _25249_/A sky130_fd_sc_hd__or2_1
X_15000_ _26443_/Q _14988_/X _14989_/X _14999_/Y vssd1 vssd1 vccd1 vccd1 _26443_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25178_ _27528_/Q _27496_/Q vssd1 vssd1 vccd1 vccd1 _25179_/B sky130_fd_sc_hd__nand2_1
X_13192_ _13192_/A vssd1 vssd1 vccd1 vccd1 _27042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24129_ _24129_/A vssd1 vssd1 vccd1 vccd1 _27338_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16951_ _24611_/A vssd1 vssd1 vccd1 vccd1 _19313_/A sky130_fd_sc_hd__buf_2
XFILLER_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15902_ _15906_/A vssd1 vssd1 vccd1 vccd1 _15902_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19670_ _19659_/X _19661_/X _19663_/X _19665_/X _19666_/X _19667_/X vssd1 vssd1 vccd1
+ vccd1 _19671_/A sky130_fd_sc_hd__mux4_1
X_16882_ _16835_/A _16599_/A _16647_/X _16881_/X vssd1 vssd1 vccd1 vccd1 _16882_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18621_ _18689_/S vssd1 vssd1 vccd1 vccd1 _18630_/S sky130_fd_sc_hd__clkbuf_2
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27819_ _25716_/X _27819_/D vssd1 vssd1 vccd1 vccd1 _27819_/Q sky130_fd_sc_hd__dfxtp_1
X_15833_ _15833_/A vssd1 vssd1 vccd1 vccd1 _26084_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _26712_/Q _26680_/Q _26648_/Q _26616_/Q _18345_/X _18012_/A vssd1 vssd1 vccd1
+ vccd1 _18553_/A sky130_fd_sc_hd__mux4_1
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15764_/A _15771_/B vssd1 vssd1 vccd1 vccd1 _15764_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _27809_/Q _12976_/B vssd1 vssd1 vccd1 vccd1 _12977_/A sky130_fd_sc_hd__and2_1
XFILLER_73_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17503_ _17503_/A vssd1 vssd1 vccd1 vccd1 _25835_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14715_/A vssd1 vssd1 vccd1 vccd1 _14715_/X sky130_fd_sc_hd__buf_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18483_ _18483_/A vssd1 vssd1 vccd1 vccd1 _18483_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15695_ _15695_/A _15695_/B _15695_/C _15695_/D vssd1 vssd1 vccd1 vccd1 _15712_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_75_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17434_ _27411_/Q vssd1 vssd1 vccd1 vccd1 _17434_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14646_ _15718_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14646_/Y sky130_fd_sc_hd__nor2_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17365_ _27095_/Q _27127_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17365_/X sky130_fd_sc_hd__mux2_1
XANTENNA_19 _25992_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ _15738_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14577_/Y sky130_fd_sc_hd__nor2_1
X_19104_ _19101_/X _19103_/X _19173_/S vssd1 vssd1 vccd1 vccd1 _19104_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16316_ _25973_/Q _16311_/X _16315_/X vssd1 vssd1 vccd1 vccd1 _16792_/B sky130_fd_sc_hd__a21oi_2
X_13528_ _13553_/A vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17296_ _17294_/X _17295_/X _17296_/S vssd1 vssd1 vccd1 vccd1 _17296_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19035_ _19290_/A vssd1 vssd1 vccd1 vccd1 _19035_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16247_ _16242_/S _16243_/Y _16244_/X _16245_/X _16246_/X vssd1 vssd1 vccd1 vccd1
+ _16460_/B sky130_fd_sc_hd__o41a_1
X_13459_ _14438_/A vssd1 vssd1 vccd1 vccd1 _13874_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16178_ _27520_/Q _27576_/Q vssd1 vssd1 vccd1 vccd1 _16178_/X sky130_fd_sc_hd__or2b_1
XFILLER_115_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _26389_/Q _13334_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15130_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19937_ _19937_/A vssd1 vssd1 vccd1 vccd1 _19937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19868_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19868_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18819_ _26266_/Q _26234_/Q _26202_/Q _26170_/Q _18816_/X _18818_/X vssd1 vssd1 vccd1
+ vccd1 _18819_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19799_ _19815_/A vssd1 vssd1 vccd1 vccd1 _19799_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21830_ _21899_/A vssd1 vssd1 vccd1 vccd1 _21830_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21761_ _22019_/A vssd1 vssd1 vccd1 vccd1 _21827_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20712_ _20703_/X _20705_/X _20707_/X _20709_/X _20710_/X _20711_/X vssd1 vssd1 vccd1
+ vccd1 _20713_/A sky130_fd_sc_hd__mux4_1
X_23500_ _27193_/Q _23500_/B vssd1 vssd1 vccd1 vccd1 _23500_/X sky130_fd_sc_hd__or2_1
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24480_ _24480_/A vssd1 vssd1 vccd1 vccd1 _24509_/B sky130_fd_sc_hd__clkbuf_2
X_21692_ _21740_/A vssd1 vssd1 vccd1 vccd1 _21692_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23431_ _17047_/S _23429_/X _23430_/X _23421_/X vssd1 vssd1 vccd1 vccd1 _27166_/D
+ sky130_fd_sc_hd__o211a_1
X_20643_ _20643_/A vssd1 vssd1 vccd1 vccd1 _20643_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26150_ _19841_/X _26150_/D vssd1 vssd1 vccd1 vccd1 _26150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23362_ _27779_/Q vssd1 vssd1 vccd1 vccd1 _24947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20574_ _20566_/X _20567_/X _20568_/X _20569_/X _20570_/X _20571_/X vssd1 vssd1 vccd1
+ vccd1 _20575_/A sky130_fd_sc_hd__mux4_1
X_22313_ _22299_/X _22300_/X _22301_/X _22302_/X _22303_/X _22304_/X vssd1 vssd1 vccd1
+ vccd1 _22314_/A sky130_fd_sc_hd__mux4_1
X_25101_ _25099_/X _25100_/X _27231_/Q vssd1 vssd1 vccd1 vccd1 _25101_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26081_ _19598_/X _26081_/D vssd1 vssd1 vccd1 vccd1 _26081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23293_ _23293_/A _23293_/B _23293_/C _23293_/D vssd1 vssd1 vccd1 vccd1 _23321_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_194_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25032_ _25075_/A vssd1 vssd1 vccd1 vccd1 _25067_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_106_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22244_ _22244_/A vssd1 vssd1 vccd1 vccd1 _22244_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22175_ _22175_/A vssd1 vssd1 vccd1 vccd1 _22175_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21126_ _21126_/A vssd1 vssd1 vccd1 vccd1 _21126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26983_ _22748_/X _26983_/D vssd1 vssd1 vccd1 vccd1 _26983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25934_ _25935_/CLK _25934_/D vssd1 vssd1 vccd1 vccd1 _25934_/Q sky130_fd_sc_hd__dfxtp_1
X_21057_ _21143_/A vssd1 vssd1 vccd1 vccd1 _21125_/A sky130_fd_sc_hd__buf_2
XFILLER_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20008_ _20266_/A vssd1 vssd1 vccd1 vccd1 _20076_/A sky130_fd_sc_hd__buf_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25865_ _25897_/CLK _25865_/D vssd1 vssd1 vccd1 vccd1 _25865_/Q sky130_fd_sc_hd__dfxtp_1
X_27604_ _27604_/CLK _27604_/D vssd1 vssd1 vccd1 vccd1 _27604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24816_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24914_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25796_ _25796_/A vssd1 vssd1 vccd1 vccd1 _27852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27535_ _27610_/CLK _27535_/D vssd1 vssd1 vccd1 vccd1 _27535_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24747_ _27613_/Q _24742_/X _24744_/Y _24746_/X vssd1 vssd1 vccd1 vccd1 _27613_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _21949_/X _21950_/X _21951_/X _21952_/X _21953_/X _21954_/X vssd1 vssd1 vccd1
+ vccd1 _21960_/A sky130_fd_sc_hd__mux4_1
XFILLER_188_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14500_/A vssd1 vssd1 vccd1 vccd1 _15758_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15549_/S sky130_fd_sc_hd__clkbuf_2
X_27466_ _27472_/CLK _27466_/D vssd1 vssd1 vccd1 vccd1 _27466_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24678_ _27588_/Q _24673_/X _24675_/X _24677_/X vssd1 vssd1 vccd1 vccd1 _27588_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _15708_/A _14446_/B vssd1 vssd1 vccd1 vccd1 _14431_/Y sky130_fd_sc_hd__nor2_1
X_26417_ _20765_/X _26417_/D vssd1 vssd1 vccd1 vccd1 _26417_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23629_ _23638_/C _23629_/B vssd1 vssd1 vccd1 vccd1 _27228_/D sky130_fd_sc_hd__nor2_1
XFILLER_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27397_ _27397_/CLK _27397_/D vssd1 vssd1 vccd1 vccd1 _27397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17150_ _27077_/Q _27109_/Q _17173_/S vssd1 vssd1 vccd1 vccd1 _17150_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14362_ _26670_/Q _14352_/X _14358_/X _14361_/Y vssd1 vssd1 vccd1 vccd1 _26670_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26348_ _20527_/X _26348_/D vssd1 vssd1 vccd1 vccd1 _26348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 la1_data_in[17] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
XFILLER_7_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16101_ _16790_/A vssd1 vssd1 vccd1 vccd1 _16308_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 la1_data_in[27] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
X_13313_ _27004_/Q _13228_/X _13313_/S vssd1 vssd1 vccd1 vccd1 _13314_/A sky130_fd_sc_hd__mux2_1
Xinput39 la1_data_in[8] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_4
X_14293_ _26695_/Q _14283_/X _14284_/X _14292_/Y vssd1 vssd1 vccd1 vccd1 _26695_/D
+ sky130_fd_sc_hd__a31o_1
X_17081_ _17291_/A vssd1 vssd1 vccd1 vccd1 _17081_/X sky130_fd_sc_hd__buf_2
XFILLER_122_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26279_ _20285_/X _26279_/D vssd1 vssd1 vccd1 vccd1 _26279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ _27265_/Q _13244_/B vssd1 vssd1 vccd1 vccd1 _13672_/B sky130_fd_sc_hd__nand2_1
X_16032_ _16233_/C vssd1 vssd1 vccd1 vccd1 _16298_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_28018_ _28018_/A _15985_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _13175_/A vssd1 vssd1 vccd1 vccd1 _27045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17983_ _17983_/A _17935_/X vssd1 vssd1 vccd1 vccd1 _17983_/X sky130_fd_sc_hd__or2b_1
X_19722_ _19710_/X _19711_/X _19712_/X _19713_/X _19714_/X _19715_/X vssd1 vssd1 vccd1
+ vccd1 _19723_/A sky130_fd_sc_hd__mux4_1
X_16934_ _24206_/A _27593_/Q _18489_/A _27488_/Q vssd1 vssd1 vccd1 vccd1 _16934_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19653_ _19653_/A vssd1 vssd1 vccd1 vccd1 _19653_/X sky130_fd_sc_hd__clkbuf_1
X_16865_ _16647_/A _16862_/Y _16863_/Y _16864_/Y _16641_/A vssd1 vssd1 vccd1 vccd1
+ _24218_/A sky130_fd_sc_hd__o32a_1
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18604_ _27753_/Q _18594_/X _25110_/B _25623_/S vssd1 vssd1 vccd1 vccd1 _18604_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15816_ _13139_/X _26091_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15817_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19584_ _19584_/A vssd1 vssd1 vccd1 vccd1 _19584_/X sky130_fd_sc_hd__clkbuf_1
X_16796_ _16796_/A _16916_/A vssd1 vssd1 vccd1 vccd1 _16800_/C sky130_fd_sc_hd__xnor2_1
X_18535_ _18535_/A _18474_/X vssd1 vssd1 vccd1 vccd1 _18535_/X sky130_fd_sc_hd__or2b_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _24980_/S vssd1 vssd1 vccd1 vccd1 _15747_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _27817_/Q _12965_/B vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__and2_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18466_ _18509_/A _18466_/B _18466_/C vssd1 vssd1 vccd1 vccd1 _18467_/A sky130_fd_sc_hd__and3_1
X_15678_ _13198_/X _26145_/Q _15678_/S vssd1 vssd1 vccd1 vccd1 _15679_/A sky130_fd_sc_hd__mux2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_291 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17417_ _27399_/Q _27398_/Q _27397_/Q _27396_/Q vssd1 vssd1 vccd1 vccd1 _17418_/C
+ sky130_fd_sc_hd__or4_1
X_14629_ _26584_/Q _14615_/X _14624_/X _14628_/Y vssd1 vssd1 vccd1 vccd1 _26584_/D
+ sky130_fd_sc_hd__a31o_1
X_18397_ _18389_/X _18391_/X _18396_/X _18285_/X _18372_/X vssd1 vssd1 vccd1 vccd1
+ _18398_/C sky130_fd_sc_hd__a221o_1
XFILLER_92_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17348_ _17348_/A vssd1 vssd1 vccd1 vccd1 _27943_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_158_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17279_ _17277_/X _17279_/B vssd1 vssd1 vccd1 vccd1 _17279_/X sky130_fd_sc_hd__and2b_1
XFILLER_174_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19018_ _26945_/Q _26913_/Q _26881_/Q _26849_/Q _18875_/X _18972_/X vssd1 vssd1 vccd1
+ vccd1 _19018_/X sky130_fd_sc_hd__mux4_2
XFILLER_173_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20290_ _20322_/A vssd1 vssd1 vccd1 vccd1 _20290_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23980_ _23978_/X _23979_/X _23987_/S vssd1 vssd1 vccd1 vccd1 _23980_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22931_ _22923_/X _22924_/X _22925_/X _22926_/X _22927_/X _22928_/X vssd1 vssd1 vccd1
+ vccd1 _22932_/A sky130_fd_sc_hd__mux4_1
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25650_ _25650_/A vssd1 vssd1 vccd1 vccd1 _25650_/X sky130_fd_sc_hd__clkbuf_1
X_22862_ _22862_/A vssd1 vssd1 vccd1 vccd1 _22862_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24601_ _27660_/Q _24609_/B vssd1 vssd1 vccd1 vccd1 _24602_/A sky130_fd_sc_hd__and2_1
XFILLER_73_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21813_ _21813_/A vssd1 vssd1 vccd1 vccd1 _21813_/X sky130_fd_sc_hd__clkbuf_2
X_25581_ _25578_/X _25579_/Y _25580_/Y _25446_/X vssd1 vssd1 vccd1 vccd1 _27777_/D
+ sky130_fd_sc_hd__a211oi_1
X_22793_ _22783_/X _22784_/X _22785_/X _22786_/X _22788_/X _22790_/X vssd1 vssd1 vccd1
+ vccd1 _22794_/A sky130_fd_sc_hd__mux4_1
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27320_ _27392_/CLK _27320_/D vssd1 vssd1 vccd1 vccd1 _27320_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21744_ _22616_/A vssd1 vssd1 vccd1 vccd1 _22089_/A sky130_fd_sc_hd__clkbuf_1
X_24532_ _24631_/A _24532_/B vssd1 vssd1 vccd1 vccd1 _24533_/A sky130_fd_sc_hd__and2_1
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27251_ _27636_/CLK _27251_/D vssd1 vssd1 vccd1 vccd1 _27251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21675_ _22021_/A vssd1 vssd1 vccd1 vccd1 _21740_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24463_ _27629_/Q _24467_/B vssd1 vssd1 vccd1 vccd1 _24464_/A sky130_fd_sc_hd__and2_1
XFILLER_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26202_ _20023_/X _26202_/D vssd1 vssd1 vccd1 vccd1 _26202_/Q sky130_fd_sc_hd__dfxtp_1
X_20626_ _20617_/X _20619_/X _20621_/X _20623_/X _20624_/X _20625_/X vssd1 vssd1 vccd1
+ vccd1 _20627_/A sky130_fd_sc_hd__mux4_1
X_23414_ _23482_/A vssd1 vssd1 vccd1 vccd1 _23429_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27182_ _27185_/CLK _27182_/D vssd1 vssd1 vccd1 vccd1 _27182_/Q sky130_fd_sc_hd__dfxtp_1
X_24394_ _24394_/A _24400_/B vssd1 vssd1 vccd1 vccd1 _24395_/A sky130_fd_sc_hd__and2_1
XFILLER_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26133_ _19777_/X _26133_/D vssd1 vssd1 vccd1 vccd1 _26133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23345_ _24893_/A vssd1 vssd1 vccd1 vccd1 _24772_/A sky130_fd_sc_hd__inv_2
X_20557_ _20557_/A vssd1 vssd1 vccd1 vccd1 _20557_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26064_ _26065_/CLK _26064_/D vssd1 vssd1 vccd1 vccd1 _26064_/Q sky130_fd_sc_hd__dfxtp_1
X_23276_ _27744_/Q vssd1 vssd1 vccd1 vccd1 _23276_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20488_ _20480_/X _20481_/X _20482_/X _20483_/X _20484_/X _20485_/X vssd1 vssd1 vccd1
+ vccd1 _20489_/A sky130_fd_sc_hd__mux4_1
XFILLER_138_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22227_ _22213_/X _22214_/X _22215_/X _22216_/X _22217_/X _22218_/X vssd1 vssd1 vccd1
+ vccd1 _22228_/A sky130_fd_sc_hd__mux4_1
XFILLER_65_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25015_ _25012_/X _25014_/X _25031_/S vssd1 vssd1 vccd1 vccd1 _25015_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22158_ _22174_/A vssd1 vssd1 vccd1 vccd1 _22158_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21109_ _21125_/A vssd1 vssd1 vccd1 vccd1 _21109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_1099 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22089_ _22089_/A vssd1 vssd1 vccd1 vccd1 _22162_/A sky130_fd_sc_hd__clkbuf_2
X_14980_ _26451_/Q _14974_/X _14976_/X _14979_/Y vssd1 vssd1 vccd1 vccd1 _26451_/D
+ sky130_fd_sc_hd__a31o_1
X_26966_ _22690_/X _26966_/D vssd1 vssd1 vccd1 vccd1 _26966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ _26814_/Q _13919_/X _13925_/X _13930_/Y vssd1 vssd1 vccd1 vccd1 _26814_/D
+ sky130_fd_sc_hd__a31o_1
X_25917_ _25917_/CLK _25917_/D vssd1 vssd1 vccd1 vccd1 _25917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26897_ _22446_/X _26897_/D vssd1 vssd1 vccd1 vccd1 _26897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16650_ _16650_/A _16650_/B vssd1 vssd1 vccd1 vccd1 _16650_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13862_ _26839_/Q _13844_/X _13855_/X _13861_/Y vssd1 vssd1 vccd1 vccd1 _26839_/D
+ sky130_fd_sc_hd__a31o_1
X_25848_ _25917_/CLK _25848_/D vssd1 vssd1 vccd1 vccd1 _25848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15601_ _15601_/A vssd1 vssd1 vccd1 vccd1 _26180_/D sky130_fd_sc_hd__clkbuf_1
X_16581_ _16795_/B vssd1 vssd1 vccd1 vccd1 _16831_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25779_ _17485_/X _27845_/Q _25779_/S vssd1 vssd1 vccd1 vccd1 _25780_/A sky130_fd_sc_hd__mux2_1
X_13793_ _13844_/A vssd1 vssd1 vccd1 vccd1 _13793_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18320_ _18311_/X _18314_/X _18319_/X _18253_/X vssd1 vssd1 vccd1 vccd1 _18333_/B
+ sky130_fd_sc_hd__a211o_1
X_27518_ _27706_/CLK _27518_/D vssd1 vssd1 vccd1 vccd1 _27518_/Q sky130_fd_sc_hd__dfxtp_1
X_15532_ _13190_/X _26210_/Q _15534_/S vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__mux2_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18251_ _18251_/A _18156_/X vssd1 vssd1 vccd1 vccd1 _18251_/X sky130_fd_sc_hd__or2b_1
XFILLER_163_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15463_/A vssd1 vssd1 vccd1 vccd1 _26241_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27449_ _27452_/CLK _27449_/D vssd1 vssd1 vccd1 vccd1 _27449_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17202_ _17202_/A vssd1 vssd1 vccd1 vccd1 _27931_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14414_ _15190_/A _14534_/B vssd1 vssd1 vccd1 vccd1 _14436_/A sky130_fd_sc_hd__nand2b_2
X_18182_ _18182_/A vssd1 vssd1 vccd1 vccd1 _18182_/X sky130_fd_sc_hd__buf_2
X_15394_ _15394_/A vssd1 vssd1 vccd1 vccd1 _26272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17133_ _17094_/X _17133_/B vssd1 vssd1 vccd1 vccd1 _17133_/X sky130_fd_sc_hd__and2b_1
X_14345_ _14398_/A vssd1 vssd1 vccd1 vccd1 _14345_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17064_ input38/X vssd1 vssd1 vccd1 vccd1 _17386_/S sky130_fd_sc_hd__clkbuf_4
X_14276_ _14363_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _27481_/Q _27268_/Q vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__or2_1
XFILLER_100_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13227_ _16191_/A vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__buf_2
XFILLER_152_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _13158_/A vssd1 vssd1 vccd1 vccd1 _27048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17966_ _26398_/Q _26366_/Q _26334_/Q _26302_/Q _17877_/X _17943_/X vssd1 vssd1 vccd1
+ vccd1 _17966_/X sky130_fd_sc_hd__mux4_1
X_13089_ _13089_/A vssd1 vssd1 vccd1 vccd1 _27060_/D sky130_fd_sc_hd__clkbuf_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater404 _27358_/CLK vssd1 vssd1 vccd1 vccd1 _27365_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater415 _27333_/CLK vssd1 vssd1 vccd1 vccd1 _27334_/CLK sky130_fd_sc_hd__clkbuf_1
X_16917_ _16077_/X _16833_/A _16916_/Y _16087_/X vssd1 vssd1 vccd1 vccd1 _16917_/X
+ sky130_fd_sc_hd__a31o_1
X_19705_ _19705_/A vssd1 vssd1 vccd1 vccd1 _19705_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater426 _25963_/CLK vssd1 vssd1 vccd1 vccd1 _26056_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17897_ _18285_/A vssd1 vssd1 vccd1 vccd1 _17897_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19636_ _19636_/A vssd1 vssd1 vccd1 vccd1 _19636_/X sky130_fd_sc_hd__clkbuf_1
X_16848_ _16091_/A _16843_/B _16847_/X vssd1 vssd1 vccd1 vccd1 _16848_/X sky130_fd_sc_hd__a21o_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19567_ _19567_/A _19567_/B _19567_/C vssd1 vssd1 vccd1 vccd1 _19568_/A sky130_fd_sc_hd__and3_1
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16779_ _16779_/A _16779_/B vssd1 vssd1 vccd1 vccd1 _16779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18518_ _17912_/X _18517_/X _17915_/X vssd1 vssd1 vccd1 vccd1 _18518_/X sky130_fd_sc_hd__o21a_1
XFILLER_179_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19498_ _27821_/Q _26582_/Q _26454_/Q _26134_/Q _18922_/X _18923_/X vssd1 vssd1 vccd1
+ vccd1 _19498_/X sky130_fd_sc_hd__mux4_1
X_18449_ _18447_/X _18448_/X _18514_/S vssd1 vssd1 vccd1 vccd1 _18449_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21460_ _21476_/A vssd1 vssd1 vccd1 vccd1 _21460_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20411_ _20427_/A vssd1 vssd1 vccd1 vccd1 _20411_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21391_ _21391_/A vssd1 vssd1 vccd1 vccd1 _21391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23130_ _27106_/Q _17702_/X _23132_/S vssd1 vssd1 vccd1 vccd1 _23131_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20342_ _20334_/X _20335_/X _20336_/X _20337_/X _20339_/X _20341_/X vssd1 vssd1 vccd1
+ vccd1 _20343_/A sky130_fd_sc_hd__mux4_1
XFILLER_161_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23061_ _23107_/S vssd1 vssd1 vccd1 vccd1 _23070_/S sky130_fd_sc_hd__clkbuf_2
X_20273_ _20337_/A vssd1 vssd1 vccd1 vccd1 _20273_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22012_ _22012_/A vssd1 vssd1 vccd1 vccd1 _22012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_510 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26820_ _22184_/X _26820_/D vssd1 vssd1 vccd1 vccd1 _26820_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_130_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26751_ _21942_/X _26751_/D vssd1 vssd1 vccd1 vccd1 _26751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23963_ _27087_/Q _27119_/Q _23986_/S vssd1 vssd1 vccd1 vccd1 _23963_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25702_ _25702_/A vssd1 vssd1 vccd1 vccd1 _25702_/X sky130_fd_sc_hd__clkbuf_1
X_22914_ _22914_/A vssd1 vssd1 vccd1 vccd1 _22914_/X sky130_fd_sc_hd__clkbuf_1
X_26682_ _21700_/X _26682_/D vssd1 vssd1 vccd1 vccd1 _26682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23894_ _27080_/Q _23860_/X _23861_/X _27112_/Q _23862_/X vssd1 vssd1 vccd1 vccd1
+ _23894_/X sky130_fd_sc_hd__a221o_1
XFILLER_112_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25633_ _23025_/X _23026_/X _23027_/X _23028_/X _23029_/X _23030_/X vssd1 vssd1 vccd1
+ vccd1 _25634_/A sky130_fd_sc_hd__mux4_1
XFILLER_140_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22845_ _22837_/X _22838_/X _22839_/X _22840_/X _22841_/X _22842_/X vssd1 vssd1 vccd1
+ vccd1 _22846_/A sky130_fd_sc_hd__mux4_1
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25564_ _25564_/A vssd1 vssd1 vccd1 vccd1 _25564_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22776_ _22776_/A vssd1 vssd1 vccd1 vccd1 _22776_/X sky130_fd_sc_hd__clkbuf_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27303_ _27357_/CLK _27303_/D vssd1 vssd1 vccd1 vccd1 _27303_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24515_ _27606_/Q _24554_/B vssd1 vssd1 vccd1 vccd1 _24516_/A sky130_fd_sc_hd__and2_1
X_21727_ _21721_/X _21722_/X _21723_/X _21724_/X _21725_/X _21726_/X vssd1 vssd1 vccd1
+ vccd1 _21728_/A sky130_fd_sc_hd__mux4_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25495_ _25487_/X _25492_/X _25493_/X _24870_/B _25494_/X vssd1 vssd1 vccd1 vccd1
+ _25495_/X sky130_fd_sc_hd__o311a_1
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27234_ _27236_/CLK _27234_/D vssd1 vssd1 vccd1 vccd1 _27234_/Q sky130_fd_sc_hd__dfxtp_1
X_21658_ _21658_/A vssd1 vssd1 vccd1 vccd1 _21658_/X sky130_fd_sc_hd__clkbuf_1
X_24446_ _24446_/A vssd1 vssd1 vccd1 vccd1 _27500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20609_ _20609_/A vssd1 vssd1 vccd1 vccd1 _20609_/X sky130_fd_sc_hd__clkbuf_1
X_27165_ _27642_/CLK _27165_/D vssd1 vssd1 vccd1 vccd1 _27165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21589_ _21580_/X _21582_/X _21584_/X _21586_/X _21587_/X _21588_/X vssd1 vssd1 vccd1
+ vccd1 _21590_/A sky130_fd_sc_hd__mux4_1
X_24377_ _24377_/A vssd1 vssd1 vccd1 vccd1 _27470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14130_ _14157_/A vssd1 vssd1 vccd1 vccd1 _14130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26116_ _19719_/X _26116_/D vssd1 vssd1 vccd1 vccd1 _26116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23328_ input71/X input72/X input42/X input43/X vssd1 vssd1 vccd1 vccd1 _23331_/B
+ sky130_fd_sc_hd__or4_1
X_27096_ _27096_/CLK _27096_/D vssd1 vssd1 vccd1 vccd1 _27096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14061_ _26778_/Q _14058_/X _13954_/B _14060_/Y vssd1 vssd1 vccd1 vccd1 _26778_/D
+ sky130_fd_sc_hd__a31o_1
X_26047_ _26047_/CLK _26047_/D vssd1 vssd1 vccd1 vccd1 _26047_/Q sky130_fd_sc_hd__dfxtp_1
X_23259_ _23254_/Y input69/X _23255_/Y input48/X _23258_/X vssd1 vssd1 vccd1 vccd1
+ _23275_/A sky130_fd_sc_hd__a221o_1
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_562 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13012_ _25106_/A vssd1 vssd1 vccd1 vccd1 _25733_/B sky130_fd_sc_hd__buf_4
X_17820_ _17779_/X _17796_/X _17817_/X _24396_/A vssd1 vssd1 vccd1 vccd1 _17858_/B
+ sky130_fd_sc_hd__a211o_1
X_27998_ _27998_/A _15883_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _25935_/Q _17750_/X _17754_/S vssd1 vssd1 vccd1 vccd1 _17752_/A sky130_fd_sc_hd__mux2_1
X_26949_ _22628_/X _26949_/D vssd1 vssd1 vccd1 vccd1 _26949_/Q sky130_fd_sc_hd__dfxtp_1
X_14963_ _26457_/Q _14957_/X _14960_/X _14962_/Y vssd1 vssd1 vccd1 vccd1 _26457_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16702_ _16852_/A _16851_/B _16395_/Y vssd1 vssd1 vccd1 vccd1 _16703_/B sky130_fd_sc_hd__o21ai_1
X_13914_ _26821_/Q _13906_/X _13912_/X _13913_/Y vssd1 vssd1 vccd1 vccd1 _26821_/D
+ sky130_fd_sc_hd__a31o_1
X_17682_ _17682_/A vssd1 vssd1 vccd1 vccd1 _25913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14894_ _14721_/X _26486_/Q _14896_/S vssd1 vssd1 vccd1 vccd1 _14895_/A sky130_fd_sc_hd__mux2_1
X_19421_ _19351_/X _19420_/X _19354_/X vssd1 vssd1 vccd1 vccd1 _19421_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16633_ _16633_/A _16815_/B vssd1 vssd1 vccd1 vccd1 _16807_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _13938_/A _13847_/B vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19352_ _19486_/A vssd1 vssd1 vccd1 vccd1 _19352_/X sky130_fd_sc_hd__clkbuf_2
X_16564_ _27400_/Q _16312_/X _16412_/X _25968_/Q _16563_/Y vssd1 vssd1 vccd1 vccd1
+ _16565_/A sky130_fd_sc_hd__a221o_1
X_13776_ _13870_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18303_ _18279_/X _18302_/X _18211_/X vssd1 vssd1 vccd1 vccd1 _18303_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15515_ _13144_/X _26218_/Q _15523_/S vssd1 vssd1 vccd1 vccd1 _15516_/A sky130_fd_sc_hd__mux2_1
XFILLER_188_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19283_ _19441_/A vssd1 vssd1 vccd1 vccd1 _19283_/X sky130_fd_sc_hd__buf_2
X_16495_ _16495_/A _16536_/B vssd1 vssd1 vccd1 vccd1 _16495_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18234_ _26537_/Q _26505_/Q _26473_/Q _27049_/Q _18233_/X _18141_/X vssd1 vssd1 vccd1
+ vccd1 _18234_/X sky130_fd_sc_hd__mux4_1
X_15446_ _15446_/A vssd1 vssd1 vccd1 vccd1 _26249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18165_ _26534_/Q _26502_/Q _26470_/Q _27046_/Q _18117_/X _18141_/X vssd1 vssd1 vccd1
+ vccd1 _18165_/X sky130_fd_sc_hd__mux4_1
X_15377_ _14769_/X _26279_/Q _15379_/S vssd1 vssd1 vccd1 vccd1 _15378_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _17116_/A vssd1 vssd1 vccd1 vccd1 _17116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14328_ _14344_/A vssd1 vssd1 vccd1 vccd1 _14412_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18096_ _17897_/X _18091_/X _18093_/X _18095_/X _17990_/X vssd1 vssd1 vccd1 vccd1
+ _18097_/C sky130_fd_sc_hd__a221o_1
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _27069_/Q _27101_/Q _17047_/S vssd1 vssd1 vccd1 vccd1 _17047_/X sky130_fd_sc_hd__mux2_1
X_14259_ _14346_/A _14263_/B vssd1 vssd1 vccd1 vccd1 _14259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18998_ _18996_/X _18997_/X _18941_/X vssd1 vssd1 vccd1 vccd1 _18998_/X sky130_fd_sc_hd__o21a_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater201 _25923_/CLK vssd1 vssd1 vccd1 vccd1 _27837_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater212 _27129_/CLK vssd1 vssd1 vccd1 vccd1 _27076_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater223 _27402_/CLK vssd1 vssd1 vccd1 vccd1 _27406_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17949_ _18481_/A vssd1 vssd1 vccd1 vccd1 _17949_/X sky130_fd_sc_hd__clkbuf_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater234 _27737_/CLK vssd1 vssd1 vccd1 vccd1 _27735_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater245 _27749_/CLK vssd1 vssd1 vccd1 vccd1 _27746_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater256 _27495_/CLK vssd1 vssd1 vccd1 vccd1 _27614_/CLK sky130_fd_sc_hd__clkbuf_1
X_20960_ _21028_/A vssd1 vssd1 vccd1 vccd1 _20960_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater267 _27174_/CLK vssd1 vssd1 vccd1 vccd1 _27593_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater278 _27531_/CLK vssd1 vssd1 vccd1 vccd1 _27610_/CLK sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater289 _27356_/CLK vssd1 vssd1 vccd1 vccd1 _27478_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_471 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19619_ _19605_/X _19606_/X _19607_/X _19608_/X _19609_/X _19610_/X vssd1 vssd1 vccd1
+ vccd1 _19620_/A sky130_fd_sc_hd__mux4_1
XFILLER_0_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20891_ _21149_/A vssd1 vssd1 vccd1 vccd1 _20956_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22630_ _22697_/A vssd1 vssd1 vccd1 vccd1 _22630_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22561_ _22609_/A vssd1 vssd1 vccd1 vccd1 _22561_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21512_ _21512_/A vssd1 vssd1 vccd1 vccd1 _21512_/X sky130_fd_sc_hd__clkbuf_1
X_24300_ _24300_/A _24302_/B vssd1 vssd1 vccd1 vccd1 _27430_/D sky130_fd_sc_hd__nor2_1
XFILLER_181_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22492_ _22508_/A vssd1 vssd1 vccd1 vccd1 _22492_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25280_ _25347_/A vssd1 vssd1 vccd1 vccd1 _25354_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21443_ _21475_/A vssd1 vssd1 vccd1 vccd1 _21443_/X sky130_fd_sc_hd__clkbuf_1
X_24231_ _24231_/A _24235_/B vssd1 vssd1 vccd1 vccd1 _27386_/D sky130_fd_sc_hd__nor2_1
XFILLER_148_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24162_ _27458_/Q _24162_/B vssd1 vssd1 vccd1 vccd1 _24163_/A sky130_fd_sc_hd__and2_1
X_21374_ _21390_/A vssd1 vssd1 vccd1 vccd1 _21374_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20325_ _20325_/A vssd1 vssd1 vccd1 vccd1 _20325_/X sky130_fd_sc_hd__clkbuf_1
X_23113_ _27098_/Q _17673_/X _23121_/S vssd1 vssd1 vccd1 vccd1 _23114_/A sky130_fd_sc_hd__mux2_1
X_24093_ _27395_/Q _24095_/B vssd1 vssd1 vccd1 vccd1 _24094_/A sky130_fd_sc_hd__and2_1
XFILLER_190_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27921_ _27921_/A _15966_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
X_23044_ _27068_/Q _17683_/X _23048_/S vssd1 vssd1 vccd1 vccd1 _23045_/A sky130_fd_sc_hd__mux2_1
X_20256_ _20248_/X _20249_/X _20250_/X _20251_/X _20253_/X _20255_/X vssd1 vssd1 vccd1
+ vccd1 _20257_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27852_ _27852_/CLK _27852_/D vssd1 vssd1 vccd1 vccd1 _27852_/Q sky130_fd_sc_hd__dfxtp_1
X_20187_ _20251_/A vssd1 vssd1 vccd1 vccd1 _20187_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26803_ _22122_/X _26803_/D vssd1 vssd1 vccd1 vccd1 _26803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27783_ _27783_/CLK _27783_/D vssd1 vssd1 vccd1 vccd1 _27783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24995_ _27068_/Q _27100_/Q _25004_/S vssd1 vssd1 vccd1 vccd1 _24995_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26734_ _21878_/X _26734_/D vssd1 vssd1 vccd1 vccd1 _26734_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23946_ _23946_/A vssd1 vssd1 vccd1 vccd1 _23946_/X sky130_fd_sc_hd__buf_2
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26665_ _21638_/X _26665_/D vssd1 vssd1 vccd1 vccd1 _26665_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23877_ _27078_/Q _27110_/Q _23892_/S vssd1 vssd1 vccd1 vccd1 _23877_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13630_ _13900_/A _13634_/B vssd1 vssd1 vccd1 vccd1 _13630_/Y sky130_fd_sc_hd__nor2_1
X_25616_ _25616_/A _25618_/B vssd1 vssd1 vccd1 vccd1 _27786_/D sky130_fd_sc_hd__nor2_1
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22828_ _22828_/A vssd1 vssd1 vccd1 vccd1 _22828_/X sky130_fd_sc_hd__clkbuf_1
X_26596_ _21400_/X _26596_/D vssd1 vssd1 vccd1 vccd1 _26596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ _13928_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13561_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25547_ _25572_/A vssd1 vssd1 vccd1 vccd1 _25547_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22759_ _22751_/X _22752_/X _22753_/X _22754_/X _22755_/X _22756_/X vssd1 vssd1 vccd1
+ vccd1 _22760_/A sky130_fd_sc_hd__mux4_1
XFILLER_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15300_ _26313_/Q _13373_/X _15306_/S vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__mux2_1
X_16280_ _16698_/A _16809_/A _16816_/A vssd1 vssd1 vccd1 vccd1 _16281_/B sky130_fd_sc_hd__or3_1
X_13492_ _27354_/Q _13450_/X _13451_/X _27322_/Q _13125_/X vssd1 vssd1 vccd1 vccd1
+ _14464_/A sky130_fd_sc_hd__a221oi_4
X_25478_ _24752_/A _25474_/X _25475_/Y _25477_/X _25467_/X vssd1 vssd1 vccd1 vccd1
+ _27760_/D sky130_fd_sc_hd__a221oi_1
XFILLER_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27217_ _27294_/CLK _27217_/D vssd1 vssd1 vccd1 vccd1 _27217_/Q sky130_fd_sc_hd__dfxtp_1
X_15231_ _15231_/A vssd1 vssd1 vccd1 vccd1 _26344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24429_ _27614_/Q _24433_/B vssd1 vssd1 vccd1 vccd1 _24430_/A sky130_fd_sc_hd__and2_1
X_27148_ _27148_/CLK _27148_/D vssd1 vssd1 vccd1 vccd1 _27148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15162_ _26374_/Q _13382_/X _15162_/S vssd1 vssd1 vccd1 vccd1 _15163_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14113_ _26760_/Q _14104_/X _14107_/X _14112_/Y vssd1 vssd1 vccd1 vccd1 _26760_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_181_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27079_ _27111_/CLK _27079_/D vssd1 vssd1 vccd1 vccd1 _27079_/Q sky130_fd_sc_hd__dfxtp_1
X_15093_ _14775_/X _26405_/Q _15101_/S vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__mux2_1
X_19970_ _19956_/X _19957_/X _19958_/X _19959_/X _19960_/X _19961_/X vssd1 vssd1 vccd1
+ vccd1 _19971_/A sky130_fd_sc_hd__mux4_1
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_464 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14044_ _14401_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14044_/Y sky130_fd_sc_hd__nor2_1
X_18921_ _26397_/Q _26365_/Q _26333_/Q _26301_/Q _18900_/X _18920_/X vssd1 vssd1 vccd1
+ vccd1 _18921_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18852_ _27794_/Q _26555_/Q _26427_/Q _26107_/Q _18793_/X _18851_/X vssd1 vssd1 vccd1
+ vccd1 _18852_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17803_ _17900_/A vssd1 vssd1 vccd1 vccd1 _18000_/A sky130_fd_sc_hd__buf_4
X_18783_ _26682_/Q _26650_/Q _26618_/Q _26586_/Q _18778_/X _18782_/X vssd1 vssd1 vccd1
+ vccd1 _18783_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15995_ _16108_/A _27539_/Q vssd1 vssd1 vccd1 vccd1 _16593_/A sky130_fd_sc_hd__nand2_1
X_17734_ _27426_/Q vssd1 vssd1 vccd1 vccd1 _17734_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14946_ _14946_/A vssd1 vssd1 vccd1 vccd1 _26463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17665_ _17514_/X _25903_/Q _17667_/S vssd1 vssd1 vccd1 vccd1 _17666_/A sky130_fd_sc_hd__mux2_1
X_14877_ _26493_/Q _13411_/X _14879_/S vssd1 vssd1 vccd1 vccd1 _14878_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_441 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16616_ _16616_/A _16616_/B vssd1 vssd1 vccd1 vccd1 _16616_/X sky130_fd_sc_hd__and2_1
XFILLER_51_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19404_ _19396_/X _19398_/X _19403_/X _19290_/X _19360_/X vssd1 vssd1 vccd1 vccd1
+ _19405_/C sky130_fd_sc_hd__a221o_1
X_13828_ _13921_/A _13838_/B vssd1 vssd1 vccd1 vccd1 _13828_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17596_ _17596_/A vssd1 vssd1 vccd1 vccd1 _25872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16547_ _16616_/B _16616_/A _16535_/B _16535_/A vssd1 vssd1 vccd1 vccd1 _16547_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_19335_ _19328_/X _19330_/X _19334_/X _19290_/X _19220_/X vssd1 vssd1 vccd1 vccd1
+ _19336_/C sky130_fd_sc_hd__a221o_1
X_13759_ _13940_/A _13759_/B vssd1 vssd1 vccd1 vccd1 _13759_/Y sky130_fd_sc_hd__nor2_1
XFILLER_189_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19266_ _19264_/X _19265_/X _19334_/S vssd1 vssd1 vccd1 vccd1 _19266_/X sky130_fd_sc_hd__mux2_1
X_16478_ _16711_/A _16411_/B _16477_/X vssd1 vssd1 vccd1 vccd1 _16719_/B sky130_fd_sc_hd__o21a_1
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _18208_/X _18212_/X _18216_/X _18168_/X _18122_/X vssd1 vssd1 vccd1 vccd1
+ _18218_/C sky130_fd_sc_hd__a221o_1
X_15429_ _26256_/Q _13350_/X _15429_/S vssd1 vssd1 vccd1 vccd1 _15430_/A sky130_fd_sc_hd__mux2_1
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19197_ _26536_/Q _26504_/Q _26472_/Q _27048_/Q _19102_/X _19148_/X vssd1 vssd1 vccd1
+ vccd1 _19197_/X sky130_fd_sc_hd__mux4_1
X_18148_ _24511_/A vssd1 vssd1 vccd1 vccd1 _18844_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18079_ _27802_/Q _26563_/Q _26435_/Q _26115_/Q _17996_/X _17997_/X vssd1 vssd1 vccd1
+ vccd1 _18079_/X sky130_fd_sc_hd__mux4_2
XFILLER_89_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20110_ _20095_/X _20097_/X _20099_/X _20101_/X _20102_/X _20103_/X vssd1 vssd1 vccd1
+ vccd1 _20111_/A sky130_fd_sc_hd__mux4_1
XFILLER_160_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21090_ _21090_/A vssd1 vssd1 vccd1 vccd1 _21090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20041_ _20041_/A vssd1 vssd1 vccd1 vccd1 _20041_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23800_ _23849_/A vssd1 vssd1 vccd1 vccd1 _23800_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_568 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24780_ _24780_/A _24786_/B vssd1 vssd1 vccd1 vccd1 _24780_/Y sky130_fd_sc_hd__nand2_1
X_21992_ _21992_/A vssd1 vssd1 vccd1 vccd1 _21992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23731_ _23731_/A vssd1 vssd1 vccd1 vccd1 _27267_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _22613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20943_ _20937_/X _20938_/X _20939_/X _20940_/X _20941_/X _20942_/X vssd1 vssd1 vccd1
+ vccd1 _20944_/A sky130_fd_sc_hd__mux4_1
XFILLER_93_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26450_ _20896_/X _26450_/D vssd1 vssd1 vccd1 vccd1 _26450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23662_ _23662_/A vssd1 vssd1 vccd1 vccd1 _27237_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20874_ _20942_/A vssd1 vssd1 vccd1 vccd1 _20874_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25401_ _25401_/A vssd1 vssd1 vccd1 vccd1 _27739_/D sky130_fd_sc_hd__clkbuf_1
X_22613_ _22613_/A vssd1 vssd1 vccd1 vccd1 _22959_/A sky130_fd_sc_hd__buf_2
X_26381_ _20645_/X _26381_/D vssd1 vssd1 vccd1 vccd1 _26381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23593_ _23593_/A vssd1 vssd1 vccd1 vccd1 _27218_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_179_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25332_ _25332_/A _27515_/Q vssd1 vssd1 vccd1 vccd1 _25332_/X sky130_fd_sc_hd__and2_1
X_22544_ _22891_/A vssd1 vssd1 vccd1 vccd1 _22611_/A sky130_fd_sc_hd__buf_2
XFILLER_50_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25263_ _25308_/A vssd1 vssd1 vccd1 vccd1 _25263_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22475_ _22507_/A vssd1 vssd1 vccd1 vccd1 _22475_/X sky130_fd_sc_hd__clkbuf_2
X_27002_ _22816_/X _27002_/D vssd1 vssd1 vccd1 vccd1 _27002_/Q sky130_fd_sc_hd__dfxtp_1
X_24214_ _24214_/A vssd1 vssd1 vccd1 vccd1 _27375_/D sky130_fd_sc_hd__clkbuf_1
X_21426_ _21426_/A vssd1 vssd1 vccd1 vccd1 _21426_/X sky130_fd_sc_hd__clkbuf_1
X_25194_ _25190_/A _25187_/X _25190_/B _25188_/A vssd1 vssd1 vccd1 vccd1 _25198_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21357_ _21389_/A vssd1 vssd1 vccd1 vccd1 _21357_/X sky130_fd_sc_hd__clkbuf_1
X_24145_ _27450_/Q _24151_/B vssd1 vssd1 vccd1 vccd1 _24146_/A sky130_fd_sc_hd__and2_1
XFILLER_146_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20308_ _20302_/X _20303_/X _20304_/X _20305_/X _20306_/X _20307_/X vssd1 vssd1 vccd1
+ vccd1 _20309_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21288_ _21304_/A vssd1 vssd1 vccd1 vccd1 _21288_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24076_ _27387_/Q _24084_/B vssd1 vssd1 vccd1 vccd1 _24077_/A sky130_fd_sc_hd__and2_1
XFILLER_146_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20239_ _20239_/A vssd1 vssd1 vccd1 vccd1 _20239_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23027_ _25637_/A vssd1 vssd1 vccd1 vccd1 _23027_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27835_ _27835_/CLK _27835_/D vssd1 vssd1 vccd1 vccd1 _27835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _14800_/A vssd1 vssd1 vccd1 vccd1 _26526_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _26107_/Q _15774_/X _15703_/B _15779_/Y vssd1 vssd1 vccd1 vccd1 _26107_/D
+ sky130_fd_sc_hd__a31o_1
X_27766_ _27766_/CLK _27766_/D vssd1 vssd1 vccd1 vccd1 _27766_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _27802_/Q _12998_/B vssd1 vssd1 vccd1 vccd1 _12993_/A sky130_fd_sc_hd__and2_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24978_ _27066_/Q _27098_/Q _25004_/S vssd1 vssd1 vccd1 vccd1 _24978_/X sky130_fd_sc_hd__mux2_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26717_ _21820_/X _26717_/D vssd1 vssd1 vccd1 vccd1 _26717_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14731_ _14731_/A vssd1 vssd1 vccd1 vccd1 _14731_/X sky130_fd_sc_hd__clkbuf_4
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23929_ _23929_/A vssd1 vssd1 vccd1 vccd1 _23929_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27697_ _27699_/CLK _27697_/D vssd1 vssd1 vccd1 vccd1 _27697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _27416_/Q vssd1 vssd1 vccd1 vccd1 _17450_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26648_ _21576_/X _26648_/D vssd1 vssd1 vccd1 vccd1 _26648_/Q sky130_fd_sc_hd__dfxtp_1
X_14662_ _15736_/A _14672_/B vssd1 vssd1 vccd1 vccd1 _14662_/Y sky130_fd_sc_hd__nor2_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _25953_/Q vssd1 vssd1 vccd1 vccd1 _16401_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ _13639_/A vssd1 vssd1 vccd1 vccd1 _13613_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17381_ _17338_/X _17381_/B vssd1 vssd1 vccd1 vccd1 _17381_/X sky130_fd_sc_hd__and2b_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14593_ _15754_/A _14597_/B vssd1 vssd1 vccd1 vccd1 _14593_/Y sky130_fd_sc_hd__nor2_1
X_26579_ _21340_/X _26579_/D vssd1 vssd1 vccd1 vccd1 _26579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19120_ _19117_/X _19119_/X _19211_/S vssd1 vssd1 vccd1 vccd1 _19120_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16332_ _16754_/A _16351_/B vssd1 vssd1 vccd1 vccd1 _16332_/X sky130_fd_sc_hd__or2_1
X_13544_ _27343_/Q _13529_/X _13530_/X _27311_/Q _13187_/X vssd1 vssd1 vccd1 vccd1
+ _14503_/A sky130_fd_sc_hd__a221oi_4
XFILLER_199_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19051_ _19123_/A _19051_/B vssd1 vssd1 vccd1 vccd1 _19051_/X sky130_fd_sc_hd__or2_1
X_16263_ _26058_/Q vssd1 vssd1 vccd1 vccd1 _16263_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13475_ _13546_/A vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_185_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18002_ _18156_/A vssd1 vssd1 vccd1 vccd1 _18580_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15214_ _15260_/S vssd1 vssd1 vccd1 vccd1 _15223_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16194_ _26045_/Q _16215_/B _16194_/C vssd1 vssd1 vccd1 vccd1 _16194_/X sky130_fd_sc_hd__and3_1
XFILLER_154_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15145_ _26382_/Q _13357_/X _15151_/S vssd1 vssd1 vccd1 vccd1 _15146_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19953_ _19953_/A vssd1 vssd1 vccd1 vccd1 _19953_/X sky130_fd_sc_hd__clkbuf_1
X_15076_ _15076_/A vssd1 vssd1 vccd1 vccd1 _26413_/D sky130_fd_sc_hd__clkbuf_1
X_14027_ _26788_/Q _14024_/X _14019_/X _14026_/Y vssd1 vssd1 vccd1 vccd1 _26788_/D
+ sky130_fd_sc_hd__a31o_1
X_18904_ _18899_/X _18902_/X _19499_/S vssd1 vssd1 vccd1 vccd1 _18904_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19884_ _19900_/A vssd1 vssd1 vccd1 vccd1 _19884_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18835_ _18827_/X _18832_/X _19539_/S vssd1 vssd1 vccd1 vccd1 _18835_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18766_ _19297_/A vssd1 vssd1 vccd1 vccd1 _19338_/A sky130_fd_sc_hd__clkbuf_2
X_15978_ _15979_/A vssd1 vssd1 vccd1 vccd1 _15978_/Y sky130_fd_sc_hd__inv_2
X_17717_ _17717_/A vssd1 vssd1 vccd1 vccd1 _25924_/D sky130_fd_sc_hd__clkbuf_1
X_14929_ _14772_/X _26470_/Q _14929_/S vssd1 vssd1 vccd1 vccd1 _14930_/A sky130_fd_sc_hd__mux2_1
X_18697_ _18697_/A vssd1 vssd1 vccd1 vccd1 _26011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17648_ _17488_/X _25895_/Q _17656_/S vssd1 vssd1 vccd1 vccd1 _17649_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17579_ _17579_/A vssd1 vssd1 vccd1 vccd1 _25864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19318_ _26702_/Q _26670_/Q _26638_/Q _26606_/Q _19317_/X _19227_/X vssd1 vssd1 vccd1
+ vccd1 _19318_/X sky130_fd_sc_hd__mux4_2
X_20590_ _20582_/X _20583_/X _20584_/X _20585_/X _20586_/X _20587_/X vssd1 vssd1 vccd1
+ vccd1 _20591_/A sky130_fd_sc_hd__mux4_2
XFILLER_32_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _26827_/Q _26795_/Q _26763_/Q _26731_/Q _19203_/X _19248_/X vssd1 vssd1 vccd1
+ vccd1 _19250_/B sky130_fd_sc_hd__mux4_2
XFILLER_31_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22260_ _22260_/A vssd1 vssd1 vccd1 vccd1 _22260_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21211_ _21211_/A vssd1 vssd1 vccd1 vccd1 _21211_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22191_ _22173_/X _22174_/X _22175_/X _22176_/X _22179_/X _22182_/X vssd1 vssd1 vccd1
+ vccd1 _22192_/A sky130_fd_sc_hd__mux4_1
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21142_ _21142_/A vssd1 vssd1 vccd1 vccd1 _21142_/X sky130_fd_sc_hd__clkbuf_2
X_21073_ _21058_/X _21060_/X _21062_/X _21064_/X _21065_/X _21066_/X vssd1 vssd1 vccd1
+ vccd1 _21074_/A sky130_fd_sc_hd__mux4_1
X_25950_ _26049_/CLK _25950_/D vssd1 vssd1 vccd1 vccd1 _25950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24901_ _27770_/Q _24902_/B vssd1 vssd1 vccd1 vccd1 _24910_/C sky130_fd_sc_hd__and2_1
X_20024_ _20009_/X _20011_/X _20013_/X _20015_/X _20016_/X _20017_/X vssd1 vssd1 vccd1
+ vccd1 _20025_/A sky130_fd_sc_hd__mux4_1
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25881_ _27135_/CLK _25881_/D vssd1 vssd1 vccd1 vccd1 _25881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27620_ _27621_/CLK _27620_/D vssd1 vssd1 vccd1 vccd1 _27620_/Q sky130_fd_sc_hd__dfxtp_1
X_24832_ _24838_/A _24832_/B vssd1 vssd1 vccd1 vccd1 _24832_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27551_ _27651_/CLK _27551_/D vssd1 vssd1 vccd1 vccd1 _27551_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24763_ _24763_/A _24772_/B vssd1 vssd1 vccd1 vccd1 _24763_/Y sky130_fd_sc_hd__nand2_1
X_21975_ _21965_/X _21966_/X _21967_/X _21968_/X _21969_/X _21970_/X vssd1 vssd1 vccd1
+ vccd1 _21976_/A sky130_fd_sc_hd__mux4_1
XFILLER_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26502_ _21072_/X _26502_/D vssd1 vssd1 vccd1 vccd1 _26502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23714_ _25601_/A _27261_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23715_/A sky130_fd_sc_hd__mux2_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20926_ _20942_/A vssd1 vssd1 vccd1 vccd1 _20926_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27482_ _27484_/CLK _27482_/D vssd1 vssd1 vccd1 vccd1 _27482_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24694_ _27179_/Q _24698_/B vssd1 vssd1 vccd1 vccd1 _24694_/X sky130_fd_sc_hd__or2_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26433_ _20829_/X _26433_/D vssd1 vssd1 vccd1 vccd1 _26433_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23645_ _23643_/X _23638_/X _23644_/Y vssd1 vssd1 vccd1 vccd1 _27231_/D sky130_fd_sc_hd__o21a_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20857_ _20857_/A vssd1 vssd1 vccd1 vccd1 _20857_/X sky130_fd_sc_hd__clkbuf_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26364_ _20581_/X _26364_/D vssd1 vssd1 vccd1 vccd1 _26364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23576_ _27772_/Q _27214_/Q _23576_/S vssd1 vssd1 vccd1 vccd1 _23577_/B sky130_fd_sc_hd__mux2_1
X_20788_ _20788_/A vssd1 vssd1 vccd1 vccd1 _22537_/A sky130_fd_sc_hd__buf_6
XFILLER_22_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25315_ _25329_/A _25329_/B _25329_/C vssd1 vssd1 vccd1 vccd1 _25319_/B sky130_fd_sc_hd__or3_1
X_22527_ _22519_/X _22520_/X _22521_/X _22522_/X _22524_/X _22526_/X vssd1 vssd1 vccd1
+ vccd1 _22528_/A sky130_fd_sc_hd__mux4_1
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26295_ _20343_/X _26295_/D vssd1 vssd1 vccd1 vccd1 _26295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25246_ _27706_/Q _25223_/X _25245_/Y _25214_/X vssd1 vssd1 vccd1 vccd1 _27706_/D
+ sky130_fd_sc_hd__o211a_1
X_13260_ _13317_/S vssd1 vssd1 vccd1 vccd1 _13269_/S sky130_fd_sc_hd__clkbuf_2
X_22458_ _22522_/A vssd1 vssd1 vccd1 vccd1 _22458_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21409_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21476_/A sky130_fd_sc_hd__clkbuf_2
X_25177_ _27528_/Q _27496_/Q vssd1 vssd1 vccd1 vccd1 _25190_/A sky130_fd_sc_hd__or2_1
X_13191_ _27042_/Q _13190_/X _13199_/S vssd1 vssd1 vccd1 vccd1 _13192_/A sky130_fd_sc_hd__mux2_1
X_22389_ _22421_/A vssd1 vssd1 vccd1 vccd1 _22389_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24128_ _27443_/Q _24128_/B vssd1 vssd1 vccd1 vccd1 _24129_/A sky130_fd_sc_hd__and2_1
XFILLER_159_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16950_ _24511_/A vssd1 vssd1 vccd1 vccd1 _24611_/A sky130_fd_sc_hd__clkbuf_4
X_24059_ _27380_/Q _24061_/B vssd1 vssd1 vccd1 vccd1 _24060_/A sky130_fd_sc_hd__and2_1
XFILLER_2_787 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15901_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15906_/A sky130_fd_sc_hd__buf_2
X_16881_ _16835_/A _16599_/A _16621_/A vssd1 vssd1 vccd1 vccd1 _16881_/X sky130_fd_sc_hd__o21ba_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18620_ _18676_/A vssd1 vssd1 vccd1 vccd1 _18689_/S sky130_fd_sc_hd__buf_2
X_15832_ _13179_/X _26084_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15833_/A sky130_fd_sc_hd__mux2_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27818_ _25714_/X _27818_/D vssd1 vssd1 vccd1 vccd1 _27818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _26840_/Q _26808_/Q _26776_/Q _26744_/Q _17832_/X _17835_/X vssd1 vssd1 vccd1
+ vccd1 _18551_/X sky130_fd_sc_hd__mux4_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _26114_/Q _15760_/X _15753_/X _15762_/Y vssd1 vssd1 vccd1 vccd1 _26114_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12975_/A vssd1 vssd1 vccd1 vccd1 _27810_/D sky130_fd_sc_hd__clkbuf_1
X_27749_ _27749_/CLK _27749_/D vssd1 vssd1 vccd1 vccd1 _27749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_569 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _17501_/X _25835_/Q _17502_/S vssd1 vssd1 vccd1 vccd1 _17503_/A sky130_fd_sc_hd__mux2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _14714_/A vssd1 vssd1 vccd1 vccd1 _26553_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _26292_/Q _26260_/Q _26228_/Q _26196_/Q _18458_/X _18481_/X vssd1 vssd1 vccd1
+ vccd1 _18482_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15694_ _15694_/A vssd1 vssd1 vccd1 vccd1 _26138_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17433_/A vssd1 vssd1 vccd1 vccd1 _25813_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ _14671_/A vssd1 vssd1 vccd1 vccd1 _14645_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17364_ _17116_/A _17359_/X _17361_/X _17363_/X vssd1 vssd1 vccd1 vccd1 _17364_/X
+ sky130_fd_sc_hd__o22a_1
X_14576_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14576_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16315_ _27405_/Q _16312_/X _16314_/X _14718_/A vssd1 vssd1 vccd1 vccd1 _16315_/X
+ sky130_fd_sc_hd__a22o_1
X_19103_ _26532_/Q _26500_/Q _26468_/Q _27044_/Q _19102_/X _19032_/X vssd1 vssd1 vccd1
+ vccd1 _19103_/X sky130_fd_sc_hd__mux4_1
X_13527_ _26950_/Q _13510_/X _13505_/X _13526_/Y vssd1 vssd1 vccd1 vccd1 _26950_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17295_ _27089_/Q _27121_/Q _17295_/S vssd1 vssd1 vccd1 vccd1 _17295_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19034_ _19031_/X _19033_/X _19057_/S vssd1 vssd1 vccd1 vccd1 _19034_/X sky130_fd_sc_hd__mux2_1
X_16246_ _27532_/Q _16034_/A vssd1 vssd1 vccd1 vccd1 _16246_/X sky130_fd_sc_hd__or2b_1
X_13458_ _27361_/Q _13450_/X _13451_/X _27329_/Q _13083_/X vssd1 vssd1 vccd1 vccd1
+ _14438_/A sky130_fd_sc_hd__a221oi_4
XFILLER_161_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16177_ _16177_/A _16191_/B _16197_/C vssd1 vssd1 vccd1 vccd1 _16177_/X sky130_fd_sc_hd__and3_1
X_13389_ _14779_/A vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15128_ _15128_/A vssd1 vssd1 vccd1 vccd1 _26390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19936_ _19918_/X _19921_/X _19924_/X _19927_/X _19928_/X _19929_/X vssd1 vssd1 vccd1
+ vccd1 _19937_/A sky130_fd_sc_hd__mux4_1
X_15059_ _15116_/S vssd1 vssd1 vccd1 vccd1 _15068_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19867_ _19899_/A vssd1 vssd1 vccd1 vccd1 _19867_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18818_ _19385_/A vssd1 vssd1 vccd1 vccd1 _18818_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19798_ _19814_/A vssd1 vssd1 vccd1 vccd1 _19798_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18749_ _26035_/Q _17756_/X _18757_/S vssd1 vssd1 vccd1 vccd1 _18750_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21760_ _21826_/A vssd1 vssd1 vccd1 vccd1 _21760_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20711_ _20759_/A vssd1 vssd1 vccd1 vccd1 _20711_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21691_ _21739_/A vssd1 vssd1 vccd1 vccd1 _21691_/X sky130_fd_sc_hd__clkbuf_1
X_23430_ _27166_/Q _23430_/B vssd1 vssd1 vccd1 vccd1 _23430_/X sky130_fd_sc_hd__or2_1
X_20642_ _20636_/X _20637_/X _20638_/X _20639_/X _20640_/X _20641_/X vssd1 vssd1 vccd1
+ vccd1 _20643_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20573_ _20573_/A vssd1 vssd1 vccd1 vccd1 _20573_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23361_ _23361_/A _23361_/B _23360_/X vssd1 vssd1 vccd1 vccd1 _23410_/A sky130_fd_sc_hd__or3b_1
XFILLER_165_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25100_ _25927_/Q _25993_/Q _25826_/Q _26025_/Q _25018_/A _25070_/X vssd1 vssd1 vccd1
+ vccd1 _25100_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22312_ _22312_/A vssd1 vssd1 vccd1 vccd1 _22312_/X sky130_fd_sc_hd__clkbuf_1
X_26080_ _19596_/X _26080_/D vssd1 vssd1 vccd1 vccd1 _26080_/Q sky130_fd_sc_hd__dfxtp_1
X_23292_ _27724_/Q _23290_/Y _23291_/Y input49/X vssd1 vssd1 vccd1 vccd1 _23293_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25031_ _25029_/X _25030_/X _25031_/S vssd1 vssd1 vccd1 vccd1 _25031_/X sky130_fd_sc_hd__mux2_2
X_22243_ _22229_/X _22230_/X _22231_/X _22232_/X _22233_/X _22234_/X vssd1 vssd1 vccd1
+ vccd1 _22244_/A sky130_fd_sc_hd__mux4_1
XFILLER_178_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22174_ _22174_/A vssd1 vssd1 vccd1 vccd1 _22174_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21125_ _21125_/A vssd1 vssd1 vccd1 vccd1 _21125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26982_ _22746_/X _26982_/D vssd1 vssd1 vccd1 vccd1 _26982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25933_ _26030_/CLK _25933_/D vssd1 vssd1 vccd1 vccd1 _25933_/Q sky130_fd_sc_hd__dfxtp_1
X_21056_ _21056_/A vssd1 vssd1 vccd1 vccd1 _21056_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20007_ _20007_/A vssd1 vssd1 vccd1 vccd1 _20007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25864_ _25897_/CLK _25864_/D vssd1 vssd1 vccd1 vccd1 _25864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27603_ _27604_/CLK _27603_/D vssd1 vssd1 vccd1 vccd1 _27603_/Q sky130_fd_sc_hd__dfxtp_1
X_24815_ _24815_/A _24815_/B vssd1 vssd1 vccd1 vccd1 _24815_/Y sky130_fd_sc_hd__nand2_1
X_25795_ _17508_/X _27852_/Q _25801_/S vssd1 vssd1 vccd1 vccd1 _25796_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27534_ _27534_/CLK _27534_/D vssd1 vssd1 vccd1 vccd1 _27534_/Q sky130_fd_sc_hd__dfxtp_2
X_24746_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24746_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21958_ _21958_/A vssd1 vssd1 vccd1 vccd1 _21958_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27465_ _27467_/CLK _27465_/D vssd1 vssd1 vccd1 vccd1 _27465_/Q sky130_fd_sc_hd__dfxtp_1
X_20909_ _20941_/A vssd1 vssd1 vccd1 vccd1 _20909_/X sky130_fd_sc_hd__clkbuf_2
X_24677_ _24729_/A vssd1 vssd1 vccd1 vccd1 _24677_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21889_ _21879_/X _21880_/X _21881_/X _21882_/X _21883_/X _21884_/X vssd1 vssd1 vccd1
+ vccd1 _21890_/A sky130_fd_sc_hd__mux4_1
XFILLER_199_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14446_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_26416_ _20763_/X _26416_/D vssd1 vssd1 vccd1 vccd1 _26416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23628_ _27227_/Q _27228_/Q _15774_/X vssd1 vssd1 vccd1 vccd1 _23629_/B sky130_fd_sc_hd__o21ai_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27396_ _27401_/CLK _27396_/D vssd1 vssd1 vccd1 vccd1 _27396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14361_/A _14363_/B vssd1 vssd1 vccd1 vccd1 _14361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26347_ _20525_/X _26347_/D vssd1 vssd1 vccd1 vccd1 _26347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23559_ _27767_/Q _27209_/Q _23559_/S vssd1 vssd1 vccd1 vccd1 _23560_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_864 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput18 la1_data_in[18] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_4
X_16100_ _27406_/Q _16094_/X _16098_/X _25974_/Q _16099_/Y vssd1 vssd1 vccd1 vccd1
+ _16790_/A sky130_fd_sc_hd__a221o_1
XFILLER_11_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13312_ _13312_/A vssd1 vssd1 vccd1 vccd1 _27005_/D sky130_fd_sc_hd__clkbuf_1
Xinput29 la1_data_in[28] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_6
X_17080_ _17080_/A vssd1 vssd1 vccd1 vccd1 _27921_/A sky130_fd_sc_hd__clkbuf_1
X_14292_ _14381_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14292_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26278_ _20283_/X _26278_/D vssd1 vssd1 vccd1 vccd1 _26278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_28017_ _28017_/A _15981_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_16031_ _16194_/C vssd1 vssd1 vccd1 vccd1 _16233_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_25229_ _25229_/A _25229_/B vssd1 vssd1 vccd1 vccd1 _25230_/B sky130_fd_sc_hd__xor2_1
X_13243_ _15334_/C _15334_/B _15045_/B vssd1 vssd1 vccd1 vccd1 _15783_/A sky130_fd_sc_hd__nand3_2
XFILLER_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13174_ _27045_/Q _13172_/X _13199_/S vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17982_ _26143_/Q _26079_/Q _27007_/Q _26975_/Q _17870_/X _17959_/X vssd1 vssd1 vccd1
+ vccd1 _17983_/A sky130_fd_sc_hd__mux4_1
XFILLER_96_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19721_ _19721_/A vssd1 vssd1 vccd1 vccd1 _19721_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16933_ _27597_/Q vssd1 vssd1 vccd1 vccd1 _18489_/A sky130_fd_sc_hd__clkinv_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19652_ _19637_/X _19638_/X _19639_/X _19640_/X _19644_/X _19647_/X vssd1 vssd1 vccd1
+ vccd1 _19653_/A sky130_fd_sc_hd__mux4_1
X_16864_ _16864_/A _16864_/B vssd1 vssd1 vccd1 vccd1 _16864_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _25625_/S vssd1 vssd1 vccd1 vccd1 _25623_/S sky130_fd_sc_hd__clkbuf_4
X_15815_ _15815_/A vssd1 vssd1 vccd1 vccd1 _26092_/D sky130_fd_sc_hd__clkbuf_1
X_16795_ _16831_/A _16795_/B vssd1 vssd1 vccd1 vccd1 _16800_/B sky130_fd_sc_hd__xnor2_1
XFILLER_93_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19583_ _19570_/X _19572_/X _19574_/X _19576_/X _19577_/X _19578_/X vssd1 vssd1 vccd1
+ vccd1 _19584_/A sky130_fd_sc_hd__mux4_1
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18534_ _26711_/Q _26679_/Q _26647_/Q _26615_/Q _18345_/X _18408_/X vssd1 vssd1 vccd1
+ vccd1 _18535_/A sky130_fd_sc_hd__mux4_1
X_15746_ _26120_/Q _15734_/X _15740_/X _15745_/Y vssd1 vssd1 vccd1 vccd1 _26120_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _12958_/A vssd1 vssd1 vccd1 vccd1 _27818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18465_ _18457_/X _18460_/X _18464_/X _18443_/X _18372_/X vssd1 vssd1 vccd1 vccd1
+ _18466_/C sky130_fd_sc_hd__a221o_1
X_15677_ _15677_/A vssd1 vssd1 vccd1 vccd1 _26146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_270 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14628_ _15701_/A _14631_/B vssd1 vssd1 vccd1 vccd1 _14628_/Y sky130_fd_sc_hd__nor2_1
X_17416_ _27395_/Q _27394_/Q _27393_/Q _27392_/Q vssd1 vssd1 vccd1 vccd1 _17418_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA_292 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18396_ _18393_/X _18394_/X _18488_/S vssd1 vssd1 vccd1 vccd1 _18396_/X sky130_fd_sc_hd__mux2_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17347_ _27222_/Q _17346_/X _17367_/S vssd1 vssd1 vccd1 vccd1 _17348_/A sky130_fd_sc_hd__mux2_1
X_14559_ _26610_/Q _14549_/X _14553_/X _14558_/Y vssd1 vssd1 vccd1 vccd1 _26610_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17278_ _25934_/Q _26000_/Q _17315_/S vssd1 vssd1 vccd1 vccd1 _17279_/B sky130_fd_sc_hd__mux2_1
XFILLER_140_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19017_ _18996_/X _19016_/X _18941_/X vssd1 vssd1 vccd1 vccd1 _19017_/X sky130_fd_sc_hd__o21a_1
X_16229_ _27384_/Q _16244_/B _16244_/C vssd1 vssd1 vccd1 vccd1 _16229_/X sky130_fd_sc_hd__and3_1
XFILLER_115_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_405 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19919_ _25655_/A vssd1 vssd1 vccd1 vccd1 _20268_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22930_ _22930_/A vssd1 vssd1 vccd1 vccd1 _22930_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22861_ _22853_/X _22854_/X _22855_/X _22856_/X _22857_/X _22858_/X vssd1 vssd1 vccd1
+ vccd1 _22862_/A sky130_fd_sc_hd__mux4_1
X_24600_ _24611_/A vssd1 vssd1 vccd1 vccd1 _24609_/B sky130_fd_sc_hd__clkbuf_1
X_21812_ _21828_/A vssd1 vssd1 vccd1 vccd1 _21812_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25580_ _25580_/A _25601_/B vssd1 vssd1 vccd1 vccd1 _25580_/Y sky130_fd_sc_hd__nor2_1
X_22792_ _22792_/A vssd1 vssd1 vccd1 vccd1 _22792_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24531_ _24554_/A _16979_/B _24545_/S vssd1 vssd1 vccd1 vccd1 _24532_/B sky130_fd_sc_hd__mux2_1
X_21743_ _21813_/A vssd1 vssd1 vccd1 vccd1 _21743_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_197_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27250_ _27250_/CLK _27250_/D vssd1 vssd1 vccd1 vccd1 _27250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24462_ _24462_/A vssd1 vssd1 vccd1 vccd1 _27507_/D sky130_fd_sc_hd__clkbuf_1
X_21674_ _22546_/A vssd1 vssd1 vccd1 vccd1 _22021_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26201_ _20021_/X _26201_/D vssd1 vssd1 vccd1 vccd1 _26201_/Q sky130_fd_sc_hd__dfxtp_1
X_23413_ _23413_/A vssd1 vssd1 vccd1 vccd1 _23482_/A sky130_fd_sc_hd__clkbuf_1
X_20625_ _20673_/A vssd1 vssd1 vccd1 vccd1 _20625_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27181_ _27185_/CLK _27181_/D vssd1 vssd1 vccd1 vccd1 _27181_/Q sky130_fd_sc_hd__dfxtp_1
X_24393_ _24393_/A vssd1 vssd1 vccd1 vccd1 _27476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26132_ _19775_/X _26132_/D vssd1 vssd1 vccd1 vccd1 _26132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23344_ _27768_/Q vssd1 vssd1 vccd1 vccd1 _24893_/A sky130_fd_sc_hd__clkbuf_4
X_20556_ _20550_/X _20551_/X _20552_/X _20553_/X _20554_/X _20555_/X vssd1 vssd1 vccd1
+ vccd1 _20557_/A sky130_fd_sc_hd__mux4_1
XFILLER_164_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26063_ _26073_/CLK _26063_/D vssd1 vssd1 vccd1 vccd1 _26063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23275_ _23275_/A _23275_/B _23275_/C _23275_/D vssd1 vssd1 vccd1 vccd1 _23322_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20487_ _20487_/A vssd1 vssd1 vccd1 vccd1 _20487_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25014_ _27070_/Q _27102_/Q _25047_/S vssd1 vssd1 vccd1 vccd1 _25014_/X sky130_fd_sc_hd__mux2_1
X_22226_ _22226_/A vssd1 vssd1 vccd1 vccd1 _22226_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22157_ _22173_/A vssd1 vssd1 vccd1 vccd1 _22157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21108_ _21108_/A vssd1 vssd1 vccd1 vccd1 _21108_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_120_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22088_ _22161_/A vssd1 vssd1 vccd1 vccd1 _22088_/X sky130_fd_sc_hd__clkbuf_2
X_26965_ _22688_/X _26965_/D vssd1 vssd1 vccd1 vccd1 _26965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ _13930_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _13930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21039_ _21039_/A vssd1 vssd1 vccd1 vccd1 _21039_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25916_ _26016_/CLK _25916_/D vssd1 vssd1 vccd1 vccd1 _25916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26896_ _22444_/X _26896_/D vssd1 vssd1 vccd1 vccd1 _26896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ _13861_/A _13861_/B vssd1 vssd1 vccd1 vccd1 _13861_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25847_ _25878_/CLK _25847_/D vssd1 vssd1 vccd1 vccd1 _25847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15600_ _26180_/Q _14779_/A _15606_/S vssd1 vssd1 vccd1 vccd1 _15601_/A sky130_fd_sc_hd__mux2_1
X_16580_ _25970_/Q _16311_/X _16579_/X vssd1 vssd1 vccd1 vccd1 _16795_/B sky130_fd_sc_hd__a21oi_2
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25778_ _25778_/A vssd1 vssd1 vccd1 vccd1 _27844_/D sky130_fd_sc_hd__clkbuf_1
X_13792_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15531_ _15531_/A vssd1 vssd1 vccd1 vccd1 _26211_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27517_ _27706_/CLK _27517_/D vssd1 vssd1 vccd1 vccd1 _27517_/Q sky130_fd_sc_hd__dfxtp_1
X_24729_ _24729_/A vssd1 vssd1 vccd1 vccd1 _24729_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _26698_/Q _26666_/Q _26634_/Q _26602_/Q _18177_/X _18249_/X vssd1 vssd1 vccd1
+ vccd1 _18251_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ _26241_/Q _13398_/X _15462_/S vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27448_ _27461_/CLK _27448_/D vssd1 vssd1 vccd1 vccd1 _27448_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _27210_/Q _17199_/X _17250_/S vssd1 vssd1 vccd1 vccd1 _17202_/A sky130_fd_sc_hd__mux2_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14413_ _26650_/Q _14405_/X _14335_/B _14412_/Y vssd1 vssd1 vccd1 vccd1 _26650_/D
+ sky130_fd_sc_hd__a31o_1
X_18181_ _18150_/X _18174_/X _18180_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _18193_/B
+ sky130_fd_sc_hd__a211o_1
X_15393_ _14791_/X _26272_/Q _15401_/S vssd1 vssd1 vccd1 vccd1 _15394_/A sky130_fd_sc_hd__mux2_1
X_27379_ _27379_/CLK _27379_/D vssd1 vssd1 vccd1 vccd1 _27379_/Q sky130_fd_sc_hd__dfxtp_2
X_17132_ _25922_/Q _25988_/Q _17132_/S vssd1 vssd1 vccd1 vccd1 _17133_/B sky130_fd_sc_hd__mux2_1
XFILLER_168_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14344_ _14344_/A vssd1 vssd1 vccd1 vccd1 _14398_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17063_ _27070_/Q _27102_/Q _17112_/S vssd1 vssd1 vccd1 vccd1 _17063_/X sky130_fd_sc_hd__mux2_1
X_14275_ _26702_/Q _14270_/X _14271_/X _14274_/Y vssd1 vssd1 vccd1 vccd1 _26702_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16014_ _27481_/Q _16014_/B vssd1 vssd1 vccd1 vccd1 _16014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13226_ _27337_/Q _13193_/A _13194_/A _27305_/Q _13225_/X vssd1 vssd1 vccd1 vccd1
+ _16191_/A sky130_fd_sc_hd__a221o_1
XFILLER_152_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _27048_/Q _13156_/X _13167_/S vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _26526_/Q _26494_/Q _26462_/Q _27038_/Q _17964_/X _17843_/X vssd1 vssd1 vccd1
+ vccd1 _17965_/X sky130_fd_sc_hd__mux4_1
X_13088_ _27060_/Q _13086_/X _13112_/S vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater405 _27312_/CLK vssd1 vssd1 vccd1 vccd1 _27358_/CLK sky130_fd_sc_hd__clkbuf_1
X_19704_ _19694_/X _19695_/X _19696_/X _19697_/X _19698_/X _19699_/X vssd1 vssd1 vccd1
+ vccd1 _19705_/A sky130_fd_sc_hd__mux4_1
Xrepeater416 _27333_/CLK vssd1 vssd1 vccd1 vccd1 _25953_/CLK sky130_fd_sc_hd__clkbuf_1
X_16916_ _16916_/A vssd1 vssd1 vccd1 vccd1 _16916_/Y sky130_fd_sc_hd__inv_2
Xrepeater427 _26059_/CLK vssd1 vssd1 vccd1 vccd1 _27326_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17896_ _17779_/X _17886_/X _17895_/X _24396_/A vssd1 vssd1 vccd1 vccd1 _17918_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_120_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19635_ _19621_/X _19622_/X _19623_/X _19624_/X _19625_/X _19626_/X vssd1 vssd1 vccd1
+ vccd1 _19636_/A sky130_fd_sc_hd__mux4_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16847_ _25909_/Q _16200_/B _16759_/B _25911_/Q vssd1 vssd1 vccd1 vccd1 _16847_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19566_ _19560_/X _19562_/X _19565_/X _18895_/A _19220_/A vssd1 vssd1 vccd1 vccd1
+ _19567_/C sky130_fd_sc_hd__a221o_1
XFILLER_168_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16778_ _16778_/A _16778_/B vssd1 vssd1 vccd1 vccd1 _16778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ _26838_/Q _26806_/Q _26774_/Q _26742_/Q _18085_/X _17913_/X vssd1 vssd1 vccd1
+ vccd1 _18517_/X sky130_fd_sc_hd__mux4_2
X_15729_ _26127_/Q _15721_/X _15727_/X _15728_/Y vssd1 vssd1 vccd1 vccd1 _26127_/D
+ sky130_fd_sc_hd__a31o_1
X_19497_ _26966_/Q _26934_/Q _26902_/Q _26870_/Q _19061_/X _18920_/X vssd1 vssd1 vccd1
+ vccd1 _19497_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18448_ _26963_/Q _26931_/Q _26899_/Q _26867_/Q _17903_/X _18000_/X vssd1 vssd1 vccd1
+ vccd1 _18448_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18379_ _18379_/A vssd1 vssd1 vccd1 vccd1 _18379_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_187_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20410_ _20426_/A vssd1 vssd1 vccd1 vccd1 _20410_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21390_ _21390_/A vssd1 vssd1 vccd1 vccd1 _21390_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20341_ _20413_/A vssd1 vssd1 vccd1 vccd1 _20341_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20272_ _20272_/A vssd1 vssd1 vccd1 vccd1 _20337_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_23060_ _23060_/A vssd1 vssd1 vccd1 vccd1 _27075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22011_ _21997_/X _21998_/X _21999_/X _22000_/X _22002_/X _22004_/X vssd1 vssd1 vccd1
+ vccd1 _22012_/A sky130_fd_sc_hd__mux4_1
XFILLER_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26750_ _21940_/X _26750_/D vssd1 vssd1 vccd1 vccd1 _26750_/Q sky130_fd_sc_hd__dfxtp_1
X_23962_ _23960_/X _23961_/X _23985_/S vssd1 vssd1 vccd1 vccd1 _23962_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25701_ _25689_/X _25690_/X _25691_/X _25692_/X _25693_/X _25694_/X vssd1 vssd1 vccd1
+ vccd1 _25702_/A sky130_fd_sc_hd__mux4_1
X_22913_ _22907_/X _22908_/X _22909_/X _22910_/X _22911_/X _22912_/X vssd1 vssd1 vccd1
+ vccd1 _22914_/A sky130_fd_sc_hd__mux4_1
XFILLER_186_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26681_ _21698_/X _26681_/D vssd1 vssd1 vccd1 vccd1 _26681_/Q sky130_fd_sc_hd__dfxtp_1
X_23893_ _23891_/X _23892_/X _23893_/S vssd1 vssd1 vccd1 vccd1 _23893_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25632_ _25632_/A vssd1 vssd1 vccd1 vccd1 _25632_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22844_ _22844_/A vssd1 vssd1 vccd1 vccd1 _22844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25563_ _24790_/A _25534_/X _25559_/Y _25562_/X _25557_/X vssd1 vssd1 vccd1 vccd1
+ _27774_/D sky130_fd_sc_hd__a221oi_1
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22775_ _22767_/X _22768_/X _22769_/X _22770_/X _22771_/X _22772_/X vssd1 vssd1 vccd1
+ vccd1 _22776_/A sky130_fd_sc_hd__mux4_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27302_ _27302_/CLK _27302_/D vssd1 vssd1 vccd1 vccd1 _27302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24514_ _24514_/A vssd1 vssd1 vccd1 vccd1 _27526_/D sky130_fd_sc_hd__clkbuf_1
X_21726_ _21726_/A vssd1 vssd1 vccd1 vccd1 _21726_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25494_ _25524_/A vssd1 vssd1 vccd1 vccd1 _25494_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27233_ _27649_/CLK _27233_/D vssd1 vssd1 vccd1 vccd1 _27233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24445_ _27621_/Q _24445_/B vssd1 vssd1 vccd1 vccd1 _24446_/A sky130_fd_sc_hd__and2_1
XFILLER_200_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21657_ _21647_/X _21648_/X _21649_/X _21650_/X _21652_/X _21654_/X vssd1 vssd1 vccd1
+ vccd1 _21658_/A sky130_fd_sc_hd__mux4_1
XFILLER_200_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20608_ _20598_/X _20599_/X _20600_/X _20601_/X _20603_/X _20605_/X vssd1 vssd1 vccd1
+ vccd1 _20609_/A sky130_fd_sc_hd__mux4_1
X_27164_ _27541_/CLK _27164_/D vssd1 vssd1 vccd1 vccd1 _27164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24376_ _27570_/Q _24380_/B vssd1 vssd1 vccd1 vccd1 _24377_/A sky130_fd_sc_hd__and2_1
X_21588_ _21636_/A vssd1 vssd1 vccd1 vccd1 _21588_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26115_ _19717_/X _26115_/D vssd1 vssd1 vccd1 vccd1 _26115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23327_ input44/X input45/X input46/X input47/X vssd1 vssd1 vccd1 vccd1 _23331_/A
+ sky130_fd_sc_hd__or4_1
X_27095_ _27095_/CLK _27095_/D vssd1 vssd1 vccd1 vccd1 _27095_/Q sky130_fd_sc_hd__dfxtp_1
X_20539_ _20587_/A vssd1 vssd1 vccd1 vccd1 _20539_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _14412_/A _14060_/B vssd1 vssd1 vccd1 vccd1 _14060_/Y sky130_fd_sc_hd__nor2_1
X_26046_ _26048_/CLK _26046_/D vssd1 vssd1 vccd1 vccd1 _26046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23258_ _23256_/Y input50/X _23257_/Y input52/X vssd1 vssd1 vccd1 vccd1 _23258_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13011_ _23650_/A vssd1 vssd1 vccd1 vccd1 _25106_/A sky130_fd_sc_hd__buf_4
X_22209_ _22194_/X _22196_/X _22198_/X _22200_/X _22201_/X _22202_/X vssd1 vssd1 vccd1
+ vccd1 _22210_/A sky130_fd_sc_hd__mux4_1
XFILLER_165_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_574 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23189_ _17431_/X _27132_/Q _23193_/S vssd1 vssd1 vccd1 vccd1 _23190_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27997_ _27997_/A _15884_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
XFILLER_181_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17750_ _27431_/Q vssd1 vssd1 vccd1 vccd1 _17750_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14962_ _15699_/A _14966_/B vssd1 vssd1 vccd1 vccd1 _14962_/Y sky130_fd_sc_hd__nor2_1
X_26948_ _22626_/X _26948_/D vssd1 vssd1 vccd1 vccd1 _26948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16701_ _16647_/X _16808_/A _16699_/Y _16700_/Y _16641_/A vssd1 vssd1 vccd1 vccd1
+ _24242_/A sky130_fd_sc_hd__o32a_1
X_13913_ _13913_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _13913_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17681_ _25913_/Q _17680_/X _17690_/S vssd1 vssd1 vccd1 vccd1 _17682_/A sky130_fd_sc_hd__mux2_1
X_14893_ _14893_/A vssd1 vssd1 vccd1 vccd1 _26487_/D sky130_fd_sc_hd__clkbuf_1
X_26879_ _22384_/X _26879_/D vssd1 vssd1 vccd1 vccd1 _26879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19420_ _26290_/Q _26258_/Q _26226_/Q _26194_/Q _19283_/X _19352_/X vssd1 vssd1 vccd1
+ vccd1 _19420_/X sky130_fd_sc_hd__mux4_1
X_13844_ _13844_/A vssd1 vssd1 vccd1 vccd1 _13844_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16632_ _16633_/A _16632_/B vssd1 vssd1 vccd1 vccd1 _16807_/B sky130_fd_sc_hd__and2_1
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27948__434 vssd1 vssd1 vccd1 vccd1 _27948__434/HI _27948_/A sky130_fd_sc_hd__conb_1
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19351_ _19485_/A vssd1 vssd1 vccd1 vccd1 _19351_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13775_ _26870_/Q _13761_/X _13764_/X _13774_/Y vssd1 vssd1 vccd1 vccd1 _26870_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16563_ _16563_/A _16563_/B vssd1 vssd1 vccd1 vccd1 _16563_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18302_ _26284_/Q _26252_/Q _26220_/Q _26188_/Q _18301_/X _18209_/X vssd1 vssd1 vccd1
+ vccd1 _18302_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15514_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15523_/S sky130_fd_sc_hd__clkbuf_2
X_16494_ _16494_/A _16494_/B vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19282_ _19419_/A _19282_/B vssd1 vssd1 vccd1 vccd1 _19282_/X sky130_fd_sc_hd__or2_1
XFILLER_71_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _26249_/Q _13373_/X _15451_/S vssd1 vssd1 vccd1 vccd1 _15446_/A sky130_fd_sc_hd__mux2_1
X_18233_ _18392_/A vssd1 vssd1 vccd1 vccd1 _18233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15376_ _15376_/A vssd1 vssd1 vccd1 vccd1 _26280_/D sky130_fd_sc_hd__clkbuf_1
X_18164_ _18162_/X _18163_/X _18070_/X vssd1 vssd1 vccd1 vccd1 _18164_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14327_ _14813_/B _14534_/B vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__nand2b_2
X_17115_ _17115_/A vssd1 vssd1 vccd1 vccd1 _27924_/A sky130_fd_sc_hd__clkbuf_1
X_18095_ _17827_/X _18094_/X _17838_/X vssd1 vssd1 vccd1 vccd1 _18095_/X sky130_fd_sc_hd__o21a_1
XFILLER_184_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17046_ _16985_/X _17040_/X _17042_/X _17045_/X vssd1 vssd1 vccd1 vccd1 _17046_/X
+ sky130_fd_sc_hd__o22a_1
X_14258_ _14311_/A vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13209_ _27340_/Q _13193_/X _13194_/X _27308_/Q _13208_/X vssd1 vssd1 vccd1 vccd1
+ _16224_/A sky130_fd_sc_hd__a221o_4
XFILLER_131_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14189_ _14215_/A vssd1 vssd1 vccd1 vccd1 _14200_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18997_ _26688_/Q _26656_/Q _26624_/Q _26592_/Q _18847_/X _18939_/X vssd1 vssd1 vccd1
+ vccd1 _18997_/X sky130_fd_sc_hd__mux4_2
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater202 _26020_/CLK vssd1 vssd1 vccd1 vccd1 _25923_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater213 _27232_/CLK vssd1 vssd1 vccd1 vccd1 _27129_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _17948_/A vssd1 vssd1 vccd1 vccd1 _25947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater224 _27332_/CLK vssd1 vssd1 vccd1 vccd1 _27402_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater235 _27737_/CLK vssd1 vssd1 vccd1 vccd1 _27748_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater246 _27747_/CLK vssd1 vssd1 vccd1 vccd1 _27749_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater257 _27612_/CLK vssd1 vssd1 vccd1 vccd1 _27495_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater268 _27174_/CLK vssd1 vssd1 vccd1 vccd1 _27597_/CLK sky130_fd_sc_hd__clkbuf_1
X_17879_ _17876_/X _17878_/X _18568_/S vssd1 vssd1 vccd1 vccd1 _17879_/X sky130_fd_sc_hd__mux2_2
Xrepeater279 _27531_/CLK vssd1 vssd1 vccd1 vccd1 _27574_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19618_ _19618_/A vssd1 vssd1 vccd1 vccd1 _19618_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_483 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20890_ _20955_/A vssd1 vssd1 vccd1 vccd1 _20890_/X sky130_fd_sc_hd__clkbuf_1
X_19549_ _19567_/A _19549_/B _19549_/C vssd1 vssd1 vccd1 vccd1 _19550_/A sky130_fd_sc_hd__and3_1
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22560_ _22560_/A vssd1 vssd1 vccd1 vccd1 _22560_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21511_ _21494_/X _21496_/X _21498_/X _21500_/X _21501_/X _21502_/X vssd1 vssd1 vccd1
+ vccd1 _21512_/A sky130_fd_sc_hd__mux4_1
XFILLER_146_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22491_ _22507_/A vssd1 vssd1 vccd1 vccd1 _22491_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24230_ _24230_/A _24235_/B vssd1 vssd1 vccd1 vccd1 _27385_/D sky130_fd_sc_hd__nor2_1
X_21442_ _21442_/A vssd1 vssd1 vccd1 vccd1 _21442_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24161_ _24161_/A vssd1 vssd1 vccd1 vccd1 _27352_/D sky130_fd_sc_hd__clkbuf_1
X_21373_ _21389_/A vssd1 vssd1 vccd1 vccd1 _21373_/X sky130_fd_sc_hd__clkbuf_1
X_23112_ _23180_/S vssd1 vssd1 vccd1 vccd1 _23121_/S sky130_fd_sc_hd__clkbuf_2
X_20324_ _20318_/X _20319_/X _20320_/X _20321_/X _20322_/X _20323_/X vssd1 vssd1 vccd1
+ vccd1 _20325_/A sky130_fd_sc_hd__mux4_1
X_24092_ _24092_/A vssd1 vssd1 vccd1 vccd1 _27321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27920_ _27920_/A _15967_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
X_23043_ _23043_/A vssd1 vssd1 vccd1 vccd1 _27067_/D sky130_fd_sc_hd__clkbuf_1
X_20255_ _20323_/A vssd1 vssd1 vccd1 vccd1 _20255_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27851_ _27851_/CLK _27851_/D vssd1 vssd1 vccd1 vccd1 _27851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20186_ _20272_/A vssd1 vssd1 vccd1 vccd1 _20251_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26802_ _22120_/X _26802_/D vssd1 vssd1 vccd1 vccd1 _26802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27782_ _27782_/CLK _27782_/D vssd1 vssd1 vccd1 vccd1 _27782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24994_ _24992_/X _24993_/X _25003_/S vssd1 vssd1 vccd1 vccd1 _24994_/X sky130_fd_sc_hd__mux2_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26733_ _21876_/X _26733_/D vssd1 vssd1 vccd1 vccd1 _26733_/Q sky130_fd_sc_hd__dfxtp_1
X_23945_ _27846_/Q _27150_/Q _25895_/Q _25863_/Q _23920_/X _23944_/X vssd1 vssd1 vccd1
+ vccd1 _23945_/X sky130_fd_sc_hd__mux4_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26664_ _21630_/X _26664_/D vssd1 vssd1 vccd1 vccd1 _26664_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23876_ _23874_/X _23875_/X _23891_/S vssd1 vssd1 vccd1 vccd1 _23876_/X sky130_fd_sc_hd__mux2_1
X_25615_ _25615_/A _25618_/B vssd1 vssd1 vccd1 vccd1 _27785_/D sky130_fd_sc_hd__nor2_1
X_22827_ _22821_/X _22822_/X _22823_/X _22824_/X _22825_/X _22826_/X vssd1 vssd1 vccd1
+ vccd1 _22828_/A sky130_fd_sc_hd__mux4_1
X_26595_ _21398_/X _26595_/D vssd1 vssd1 vccd1 vccd1 _26595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _14515_/A vssd1 vssd1 vccd1 vccd1 _13928_/A sky130_fd_sc_hd__buf_2
X_25546_ _27708_/Q _25539_/X _25540_/X vssd1 vssd1 vccd1 vccd1 _25546_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22758_ _22758_/A vssd1 vssd1 vccd1 vccd1 _22758_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21709_ _21725_/A vssd1 vssd1 vccd1 vccd1 _21709_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _26958_/Q _13487_/X _13482_/X _13490_/Y vssd1 vssd1 vccd1 vccd1 _26958_/D
+ sky130_fd_sc_hd__a31o_1
X_25477_ _25470_/X _25166_/B _25476_/X _25452_/X vssd1 vssd1 vccd1 vccd1 _25477_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22689_ _22681_/X _22682_/X _22683_/X _22684_/X _22685_/X _22686_/X vssd1 vssd1 vccd1
+ vccd1 _22690_/A sky130_fd_sc_hd__mux4_1
XFILLER_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15230_ _14766_/X _26344_/Q _15234_/S vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27216_ _27219_/CLK _27216_/D vssd1 vssd1 vccd1 vccd1 _27216_/Q sky130_fd_sc_hd__dfxtp_1
X_24428_ _24428_/A vssd1 vssd1 vccd1 vccd1 _27492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_463 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27147_ _27845_/CLK _27147_/D vssd1 vssd1 vccd1 vccd1 _27147_/Q sky130_fd_sc_hd__dfxtp_1
X_15161_ _15161_/A vssd1 vssd1 vccd1 vccd1 _26375_/D sky130_fd_sc_hd__clkbuf_1
X_24359_ _27562_/Q _24361_/B vssd1 vssd1 vccd1 vccd1 _24360_/A sky130_fd_sc_hd__and2_1
XFILLER_138_485 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14112_ _14376_/A _14112_/B vssd1 vssd1 vccd1 vccd1 _14112_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27078_ _27111_/CLK _27078_/D vssd1 vssd1 vccd1 vccd1 _27078_/Q sky130_fd_sc_hd__dfxtp_1
X_15092_ _15103_/A vssd1 vssd1 vccd1 vccd1 _15101_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_158_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26029_ _27122_/CLK _26029_/D vssd1 vssd1 vccd1 vccd1 _26029_/Q sky130_fd_sc_hd__dfxtp_1
X_14043_ _14515_/A vssd1 vssd1 vccd1 vccd1 _14401_/A sky130_fd_sc_hd__clkbuf_2
X_18920_ _19445_/A vssd1 vssd1 vccd1 vccd1 _18920_/X sky130_fd_sc_hd__buf_6
XFILLER_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18851_ _19321_/A vssd1 vssd1 vccd1 vccd1 _18851_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17802_ _27594_/Q vssd1 vssd1 vccd1 vccd1 _17900_/A sky130_fd_sc_hd__clkbuf_2
X_18782_ _19227_/A vssd1 vssd1 vccd1 vccd1 _18782_/X sky130_fd_sc_hd__buf_4
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15994_ _16242_/S vssd1 vssd1 vccd1 vccd1 _16108_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17733_ _17733_/A vssd1 vssd1 vccd1 vccd1 _25929_/D sky130_fd_sc_hd__clkbuf_1
X_14945_ _14795_/X _26463_/Q _14951_/S vssd1 vssd1 vccd1 vccd1 _14946_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17664_ _17664_/A vssd1 vssd1 vccd1 vccd1 _25902_/D sky130_fd_sc_hd__clkbuf_1
X_14876_ _14876_/A vssd1 vssd1 vccd1 vccd1 _26494_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19403_ _19400_/X _19402_/X _19468_/S vssd1 vssd1 vccd1 vccd1 _19403_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16615_ _16700_/A _16514_/X _16546_/X vssd1 vssd1 vccd1 vccd1 _16885_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13827_ _13827_/A vssd1 vssd1 vccd1 vccd1 _13838_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17595_ _17517_/X _25872_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17596_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19334_ _19332_/X _19333_/X _19334_/S vssd1 vssd1 vccd1 vccd1 _19334_/X sky130_fd_sc_hd__mux2_1
X_13758_ _26875_/Q _13750_/X _13683_/B _13757_/Y vssd1 vssd1 vccd1 vccd1 _26875_/D
+ sky130_fd_sc_hd__a31o_1
X_16546_ _16631_/A _16664_/A _16543_/X _16544_/X _16545_/X vssd1 vssd1 vccd1 vccd1
+ _16546_/X sky130_fd_sc_hd__a311o_1
XFILLER_189_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19265_ _26539_/Q _26507_/Q _26475_/Q _27051_/Q _19242_/X _19148_/X vssd1 vssd1 vccd1
+ vccd1 _19265_/X sky130_fd_sc_hd__mux4_1
X_13689_ _13870_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13689_/Y sky130_fd_sc_hd__nor2_1
X_16477_ _16711_/A _16411_/B _16708_/A _16708_/B vssd1 vssd1 vccd1 vccd1 _16477_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18216_ _18213_/X _18215_/X _18216_/S vssd1 vssd1 vccd1 vccd1 _18216_/X sky130_fd_sc_hd__mux2_2
X_15428_ _15428_/A vssd1 vssd1 vccd1 vccd1 _26257_/D sky130_fd_sc_hd__clkbuf_1
X_19196_ _26408_/Q _26376_/Q _26344_/Q _26312_/Q _19170_/X _19100_/X vssd1 vssd1 vccd1
+ vccd1 _19196_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15359_ _15405_/S vssd1 vssd1 vccd1 vccd1 _15368_/S sky130_fd_sc_hd__clkbuf_2
X_18147_ _18147_/A vssd1 vssd1 vccd1 vccd1 _25955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18078_ _18078_/A vssd1 vssd1 vccd1 vccd1 _25952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17029_ _17303_/A vssd1 vssd1 vccd1 vccd1 _17029_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20040_ _20028_/X _20029_/X _20030_/X _20031_/X _20032_/X _20033_/X vssd1 vssd1 vccd1
+ vccd1 _20041_/A sky130_fd_sc_hd__mux4_1
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21991_ _21981_/X _21982_/X _21983_/X _21984_/X _21985_/X _21986_/X vssd1 vssd1 vccd1
+ vccd1 _21992_/A sky130_fd_sc_hd__mux4_1
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23730_ _27371_/Q _24050_/B vssd1 vssd1 vccd1 vccd1 _23731_/A sky130_fd_sc_hd__and2_1
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _20942_/A vssd1 vssd1 vccd1 vccd1 _20942_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_420 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23661_ _24835_/A _27237_/Q _23661_/S vssd1 vssd1 vccd1 vccd1 _23662_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20873_ _21217_/A vssd1 vssd1 vccd1 vccd1 _20942_/A sky130_fd_sc_hd__clkbuf_4
X_25400_ _27739_/Q input50/X _25402_/S vssd1 vssd1 vccd1 vccd1 _25401_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22612_ _22612_/A vssd1 vssd1 vccd1 vccd1 _22612_/X sky130_fd_sc_hd__clkbuf_1
X_26380_ _20643_/X _26380_/D vssd1 vssd1 vccd1 vccd1 _26380_/Q sky130_fd_sc_hd__dfxtp_1
X_23592_ _23596_/A _23592_/B vssd1 vssd1 vccd1 vccd1 _23593_/A sky130_fd_sc_hd__and2_1
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25331_ _25332_/A _27515_/Q vssd1 vssd1 vccd1 vccd1 _25331_/Y sky130_fd_sc_hd__nor2_1
X_22543_ _22543_/A vssd1 vssd1 vccd1 vccd1 _22891_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25262_ _27708_/Q _25223_/X _25261_/Y _25254_/X vssd1 vssd1 vccd1 vccd1 _27708_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22474_ _22522_/A vssd1 vssd1 vccd1 vccd1 _22474_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27001_ _22814_/X _27001_/D vssd1 vssd1 vccd1 vccd1 _27001_/Q sky130_fd_sc_hd__dfxtp_1
X_24213_ _27573_/Q _24233_/B vssd1 vssd1 vccd1 vccd1 _24214_/A sky130_fd_sc_hd__and2_1
XFILLER_194_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21425_ _21408_/X _21410_/X _21412_/X _21414_/X _21415_/X _21416_/X vssd1 vssd1 vccd1
+ vccd1 _21426_/A sky130_fd_sc_hd__mux4_1
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25193_ _27699_/Q _25184_/X _25192_/Y _25175_/X vssd1 vssd1 vccd1 vccd1 _27699_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24144_ _24144_/A vssd1 vssd1 vccd1 vccd1 _27344_/D sky130_fd_sc_hd__clkbuf_1
X_21356_ _21356_/A vssd1 vssd1 vccd1 vccd1 _21356_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_903 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20307_ _20323_/A vssd1 vssd1 vccd1 vccd1 _20307_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24075_ _24119_/A vssd1 vssd1 vccd1 vccd1 _24084_/B sky130_fd_sc_hd__clkbuf_1
X_21287_ _21303_/A vssd1 vssd1 vccd1 vccd1 _21287_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_542 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23026_ _25636_/A vssd1 vssd1 vccd1 vccd1 _23026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20238_ _20232_/X _20233_/X _20234_/X _20235_/X _20236_/X _20237_/X vssd1 vssd1 vccd1
+ vccd1 _20239_/A sky130_fd_sc_hd__mux4_1
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27834_ _27835_/CLK _27834_/D vssd1 vssd1 vccd1 vccd1 _27834_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ _20237_/A vssd1 vssd1 vccd1 vccd1 _20169_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12991_/A vssd1 vssd1 vccd1 vccd1 _27803_/D sky130_fd_sc_hd__clkbuf_1
X_27765_ _27768_/CLK _27765_/D vssd1 vssd1 vccd1 vccd1 _27765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24977_ _24973_/X _24976_/X _25003_/S vssd1 vssd1 vccd1 vccd1 _24977_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26716_ _21818_/X _26716_/D vssd1 vssd1 vccd1 vccd1 _26716_/Q sky130_fd_sc_hd__dfxtp_1
X_14730_ _14730_/A vssd1 vssd1 vccd1 vccd1 _26548_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23928_ _27844_/Q _27148_/Q _25893_/Q _25861_/Q _23920_/X _23897_/X vssd1 vssd1 vccd1
+ vccd1 _23928_/X sky130_fd_sc_hd__mux4_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27696_ _27699_/CLK _27696_/D vssd1 vssd1 vccd1 vccd1 _27696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14688_/A vssd1 vssd1 vccd1 vccd1 _14672_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26647_ _21574_/X _26647_/D vssd1 vssd1 vccd1 vccd1 _26647_/Q sky130_fd_sc_hd__dfxtp_1
X_23859_ _23855_/X _23857_/X _23893_/S vssd1 vssd1 vccd1 vccd1 _23859_/X sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _26929_/Q _13599_/X _13603_/X _13611_/Y vssd1 vssd1 vccd1 vccd1 _26929_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16400_ _16400_/A vssd1 vssd1 vccd1 vccd1 _16563_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17380_ _25943_/Q _26009_/Q _17380_/S vssd1 vssd1 vccd1 vccd1 _17381_/B sky130_fd_sc_hd__mux2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26578_ _21338_/X _26578_/D vssd1 vssd1 vccd1 vccd1 _26578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13543_ _26947_/Q _13535_/X _13528_/X _13542_/Y vssd1 vssd1 vccd1 vccd1 _26947_/D
+ sky130_fd_sc_hd__a31o_1
X_16331_ _16752_/A _16331_/B vssd1 vssd1 vccd1 vccd1 _16351_/B sky130_fd_sc_hd__xnor2_1
X_25529_ _27705_/Q _25509_/X _25510_/X vssd1 vssd1 vccd1 vccd1 _25529_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_30 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16262_ _16036_/X _16259_/Y _16260_/X _16261_/X vssd1 vssd1 vccd1 vccd1 _16633_/A
+ sky130_fd_sc_hd__o31a_1
X_19050_ _26146_/Q _26082_/Q _27010_/Q _26978_/Q _19049_/X _18950_/X vssd1 vssd1 vccd1
+ vccd1 _19051_/B sky130_fd_sc_hd__mux4_1
X_13474_ _14448_/A vssd1 vssd1 vccd1 vccd1 _13882_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18001_ _26944_/Q _26912_/Q _26880_/Q _26848_/Q _17999_/X _18000_/X vssd1 vssd1 vccd1
+ vccd1 _18001_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15213_ _15213_/A vssd1 vssd1 vccd1 vccd1 _26352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16193_ _16172_/X _16188_/X _16190_/Y _16191_/X _16192_/X vssd1 vssd1 vccd1 vccd1
+ _16756_/A sky130_fd_sc_hd__o41a_1
XFILLER_138_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15144_ _15144_/A vssd1 vssd1 vccd1 vccd1 _26383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19952_ _19940_/X _19941_/X _19942_/X _19943_/X _19944_/X _19945_/X vssd1 vssd1 vccd1
+ vccd1 _19953_/A sky130_fd_sc_hd__mux4_1
X_15075_ _14750_/X _26413_/Q _15079_/S vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__mux2_1
X_27991__457 vssd1 vssd1 vccd1 vccd1 _27991__457/HI _27991_/A sky130_fd_sc_hd__conb_1
X_14026_ _14388_/A _14029_/B vssd1 vssd1 vccd1 vccd1 _14026_/Y sky130_fd_sc_hd__nor2_1
X_18903_ _19296_/S vssd1 vssd1 vccd1 vccd1 _19499_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_68_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19883_ _19899_/A vssd1 vssd1 vccd1 vccd1 _19883_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18834_ _19391_/A vssd1 vssd1 vccd1 vccd1 _19539_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_110_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_490 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18765_ _18828_/A vssd1 vssd1 vccd1 vccd1 _19297_/A sky130_fd_sc_hd__buf_2
X_15977_ _15979_/A vssd1 vssd1 vccd1 vccd1 _15977_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17716_ _25924_/Q _17715_/X _17722_/S vssd1 vssd1 vccd1 vccd1 _17717_/A sky130_fd_sc_hd__mux2_1
X_14928_ _14928_/A vssd1 vssd1 vccd1 vccd1 _26471_/D sky130_fd_sc_hd__clkbuf_1
X_18696_ _26011_/Q _17680_/X _18702_/S vssd1 vssd1 vccd1 vccd1 _18697_/A sky130_fd_sc_hd__mux2_1
X_17647_ _17658_/A vssd1 vssd1 vccd1 vccd1 _17656_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14859_ _14870_/A vssd1 vssd1 vccd1 vccd1 _14868_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17578_ _17492_/X _25864_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17579_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19317_ _19317_/A vssd1 vssd1 vccd1 vccd1 _19317_/X sky130_fd_sc_hd__buf_2
XFILLER_17_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16529_ _27397_/Q _16557_/B vssd1 vssd1 vccd1 vccd1 _16529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19248_ _19407_/A vssd1 vssd1 vccd1 vccd1 _19248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19179_ _19317_/A vssd1 vssd1 vccd1 vccd1 _19179_/X sky130_fd_sc_hd__buf_2
XFILLER_157_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21210_ _21210_/A vssd1 vssd1 vccd1 vccd1 _21210_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22190_ _22190_/A vssd1 vssd1 vccd1 vccd1 _22190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21141_ _21125_/X _21126_/X _21127_/X _21128_/X _21130_/X _21132_/X vssd1 vssd1 vccd1
+ vccd1 _21142_/A sky130_fd_sc_hd__mux4_1
XFILLER_28_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21072_ _21072_/A vssd1 vssd1 vccd1 vccd1 _21072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24900_ _27656_/Q _24885_/X _24899_/Y _24890_/X vssd1 vssd1 vccd1 vccd1 _27656_/D
+ sky130_fd_sc_hd__o211a_1
X_20023_ _20023_/A vssd1 vssd1 vccd1 vccd1 _20023_/X sky130_fd_sc_hd__clkbuf_1
X_25880_ _25917_/CLK _25880_/D vssd1 vssd1 vccd1 vccd1 _25880_/Q sky130_fd_sc_hd__dfxtp_1
X_24831_ _24835_/B _24831_/B vssd1 vssd1 vccd1 vccd1 _24832_/B sky130_fd_sc_hd__xnor2_1
XFILLER_6_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24762_ _24803_/A vssd1 vssd1 vccd1 vccd1 _24772_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_27550_ _27651_/CLK _27550_/D vssd1 vssd1 vccd1 vccd1 _27550_/Q sky130_fd_sc_hd__dfxtp_1
X_21974_ _21974_/A vssd1 vssd1 vccd1 vccd1 _21974_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23713_ _23713_/A vssd1 vssd1 vccd1 vccd1 _27260_/D sky130_fd_sc_hd__clkbuf_1
X_26501_ _21070_/X _26501_/D vssd1 vssd1 vccd1 vccd1 _26501_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20925_ _20941_/A vssd1 vssd1 vccd1 vccd1 _20925_/X sky130_fd_sc_hd__clkbuf_2
X_27481_ _27520_/CLK _27481_/D vssd1 vssd1 vccd1 vccd1 _27481_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24693_ _24388_/A _24687_/X _24692_/X _24690_/X vssd1 vssd1 vccd1 vccd1 _27594_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26432_ _20827_/X _26432_/D vssd1 vssd1 vccd1 vccd1 _26432_/Q sky130_fd_sc_hd__dfxtp_1
X_23644_ _23643_/X _23638_/X _25430_/B vssd1 vssd1 vccd1 vccd1 _23644_/Y sky130_fd_sc_hd__a21oi_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20856_ _20848_/X _20849_/X _20850_/X _20851_/X _20852_/X _20853_/X vssd1 vssd1 vccd1
+ vccd1 _20857_/A sky130_fd_sc_hd__mux4_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26363_ _20579_/X _26363_/D vssd1 vssd1 vccd1 vccd1 _26363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23575_ _23575_/A vssd1 vssd1 vccd1 vccd1 _27213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20787_ _20787_/A vssd1 vssd1 vccd1 vccd1 _20787_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25314_ _27714_/Q _25308_/X _25313_/Y _25297_/X vssd1 vssd1 vccd1 vccd1 _27714_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22526_ _22598_/A vssd1 vssd1 vccd1 vccd1 _22526_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_28005__471 vssd1 vssd1 vccd1 vccd1 _28005__471/HI _28005_/A sky130_fd_sc_hd__conb_1
XFILLER_183_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26294_ _20333_/X _26294_/D vssd1 vssd1 vccd1 vccd1 _26294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25245_ _25261_/A _25245_/B vssd1 vssd1 vccd1 vccd1 _25245_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22457_ _22457_/A vssd1 vssd1 vccd1 vccd1 _22522_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21408_ _21475_/A vssd1 vssd1 vccd1 vccd1 _21408_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13190_ _14785_/A vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__buf_2
X_25176_ _27697_/Q _25142_/X _25174_/Y _25175_/X vssd1 vssd1 vccd1 vccd1 _27697_/D
+ sky130_fd_sc_hd__o211a_1
X_22388_ _22436_/A vssd1 vssd1 vccd1 vccd1 _22388_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_403 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24127_ _24127_/A vssd1 vssd1 vccd1 vccd1 _27337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21339_ _21322_/X _21324_/X _21326_/X _21328_/X _21329_/X _21330_/X vssd1 vssd1 vccd1
+ vccd1 _21340_/A sky130_fd_sc_hd__mux4_1
XFILLER_151_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24058_ _24058_/A vssd1 vssd1 vccd1 vccd1 _27306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_799 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15900_ input1/X vssd1 vssd1 vccd1 vccd1 _15925_/A sky130_fd_sc_hd__buf_2
X_23009_ _25635_/A vssd1 vssd1 vccd1 vccd1 _23009_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _16879_/A _16879_/B _16879_/C vssd1 vssd1 vccd1 vccd1 _16880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_131_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _15831_/A vssd1 vssd1 vccd1 vccd1 _26085_/D sky130_fd_sc_hd__clkbuf_1
X_27817_ _25712_/X _27817_/D vssd1 vssd1 vccd1 vccd1 _27817_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18550_ _18548_/X _18549_/X _18568_/S vssd1 vssd1 vccd1 vccd1 _18550_/X sky130_fd_sc_hd__mux2_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _15762_/A _15771_/B vssd1 vssd1 vccd1 vccd1 _15762_/Y sky130_fd_sc_hd__nor2_1
X_12974_ _27810_/Q _12976_/B vssd1 vssd1 vccd1 vccd1 _12975_/A sky130_fd_sc_hd__and2_1
X_27748_ _27748_/CLK _27748_/D vssd1 vssd1 vccd1 vccd1 _27748_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _27432_/Q vssd1 vssd1 vccd1 vccd1 _17501_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14713_ _14709_/X _26553_/Q _14725_/S vssd1 vssd1 vccd1 vccd1 _14714_/A sky130_fd_sc_hd__mux2_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18481_ _18481_/A vssd1 vssd1 vccd1 vccd1 _18481_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27679_ _27684_/CLK _27679_/D vssd1 vssd1 vccd1 vccd1 _27970_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15693_ _13240_/X _26138_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15694_/A sky130_fd_sc_hd__mux2_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17432_ _17431_/X _25813_/Q _17438_/S vssd1 vssd1 vccd1 vccd1 _17433_/A sky130_fd_sc_hd__mux2_1
X_14644_ _26579_/Q _14630_/X _14640_/X _14643_/Y vssd1 vssd1 vccd1 vccd1 _26579_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14575_ _26604_/Q _14563_/X _14566_/X _14574_/Y vssd1 vssd1 vccd1 vccd1 _26604_/D
+ sky130_fd_sc_hd__a31o_1
X_17363_ _16992_/X _17362_/X _17342_/X vssd1 vssd1 vccd1 vccd1 _17363_/X sky130_fd_sc_hd__a21bo_1
XFILLER_13_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19102_ _19414_/A vssd1 vssd1 vccd1 vccd1 _19102_/X sky130_fd_sc_hd__buf_2
XFILLER_186_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16314_ _16384_/A vssd1 vssd1 vccd1 vccd1 _16314_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13526_ _13910_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17294_ _17238_/X _17288_/X _17290_/X _17293_/X vssd1 vssd1 vccd1 vccd1 _17294_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19033_ _26529_/Q _26497_/Q _26465_/Q _27041_/Q _18984_/X _19032_/X vssd1 vssd1 vccd1
+ vccd1 _19033_/X sky130_fd_sc_hd__mux4_1
X_13457_ _13553_/A vssd1 vssd1 vccd1 vccd1 _13457_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16245_ _26055_/Q _16252_/B _16274_/C vssd1 vssd1 vccd1 vccd1 _16245_/X sky130_fd_sc_hd__and3_1
XFILLER_173_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13388_ _13388_/A vssd1 vssd1 vccd1 vccd1 _26981_/D sky130_fd_sc_hd__clkbuf_1
X_16176_ _16342_/A _16224_/B vssd1 vssd1 vccd1 vccd1 _16176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127_ _26390_/Q _13331_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15128_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19935_ _19935_/A vssd1 vssd1 vccd1 vccd1 _19935_/X sky130_fd_sc_hd__clkbuf_1
X_15058_ _15058_/A vssd1 vssd1 vccd1 vccd1 _26421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14009_ _14482_/A vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__clkbuf_2
X_19866_ _19898_/A vssd1 vssd1 vccd1 vccd1 _19866_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18817_ _18923_/A vssd1 vssd1 vccd1 vccd1 _19385_/A sky130_fd_sc_hd__buf_4
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19797_ _19813_/A vssd1 vssd1 vccd1 vccd1 _19797_/X sky130_fd_sc_hd__clkbuf_1
X_18748_ _18748_/A vssd1 vssd1 vccd1 vccd1 _18757_/S sky130_fd_sc_hd__buf_2
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18679_ _26004_/Q _17760_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _18680_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20710_ _20758_/A vssd1 vssd1 vccd1 vccd1 _20710_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21690_ _21738_/A vssd1 vssd1 vccd1 vccd1 _21690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20641_ _20673_/A vssd1 vssd1 vccd1 vccd1 _20641_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23360_ _23360_/A _23360_/B _23360_/C vssd1 vssd1 vccd1 vccd1 _23360_/X sky130_fd_sc_hd__and3_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20572_ _20566_/X _20567_/X _20568_/X _20569_/X _20570_/X _20571_/X vssd1 vssd1 vccd1
+ vccd1 _20573_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22311_ _22299_/X _22300_/X _22301_/X _22302_/X _22303_/X _22304_/X vssd1 vssd1 vccd1
+ vccd1 _22312_/A sky130_fd_sc_hd__mux4_1
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23291_ _27738_/Q vssd1 vssd1 vccd1 vccd1 _23291_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25030_ _27072_/Q _27104_/Q _25047_/S vssd1 vssd1 vccd1 vccd1 _25030_/X sky130_fd_sc_hd__mux2_1
X_22242_ _22242_/A vssd1 vssd1 vccd1 vccd1 _22242_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22173_ _22173_/A vssd1 vssd1 vccd1 vccd1 _22173_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21124_ _21124_/A vssd1 vssd1 vccd1 vccd1 _21124_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_458 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26981_ _22744_/X _26981_/D vssd1 vssd1 vccd1 vccd1 _26981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25932_ _27123_/CLK _25932_/D vssd1 vssd1 vccd1 vccd1 _25932_/Q sky130_fd_sc_hd__dfxtp_1
X_21055_ _21039_/X _21040_/X _21041_/X _21042_/X _21044_/X _21046_/X vssd1 vssd1 vccd1
+ vccd1 _21056_/A sky130_fd_sc_hd__mux4_1
XFILLER_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20006_ _19988_/X _19989_/X _19990_/X _19991_/X _19994_/X _19997_/X vssd1 vssd1 vccd1
+ vccd1 _20007_/A sky130_fd_sc_hd__mux4_1
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25863_ _25895_/CLK _25863_/D vssd1 vssd1 vccd1 vccd1 _25863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27602_ _27602_/CLK _27602_/D vssd1 vssd1 vccd1 vccd1 _27602_/Q sky130_fd_sc_hd__dfxtp_4
X_24814_ _24965_/A vssd1 vssd1 vccd1 vccd1 _24815_/A sky130_fd_sc_hd__inv_2
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25794_ _25794_/A vssd1 vssd1 vccd1 vccd1 _27851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27533_ _27539_/CLK _27533_/D vssd1 vssd1 vccd1 vccd1 _27533_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21957_ _21949_/X _21950_/X _21951_/X _21952_/X _21953_/X _21954_/X vssd1 vssd1 vccd1
+ vccd1 _21958_/A sky130_fd_sc_hd__mux4_1
X_24745_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24801_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _20956_/A vssd1 vssd1 vccd1 vccd1 _20908_/X sky130_fd_sc_hd__clkbuf_1
X_24676_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24729_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27464_ _27467_/CLK _27464_/D vssd1 vssd1 vccd1 vccd1 _27464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21888_ _21888_/A vssd1 vssd1 vccd1 vccd1 _21888_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23627_ _27227_/Q _27228_/Q vssd1 vssd1 vccd1 vccd1 _23638_/C sky130_fd_sc_hd__and2_1
X_26415_ _20761_/X _26415_/D vssd1 vssd1 vccd1 vccd1 _26415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20839_ _20839_/A vssd1 vssd1 vccd1 vccd1 _20839_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27395_ _27398_/CLK _27395_/D vssd1 vssd1 vccd1 vccd1 _27395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14360_ _26671_/Q _14352_/X _14358_/X _14359_/Y vssd1 vssd1 vccd1 vccd1 _26671_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_168_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26346_ _20523_/X _26346_/D vssd1 vssd1 vccd1 vccd1 _26346_/Q sky130_fd_sc_hd__dfxtp_1
X_23558_ _23558_/A vssd1 vssd1 vccd1 vccd1 _27208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _27005_/Q _13222_/X _13313_/S vssd1 vssd1 vccd1 vccd1 _13312_/A sky130_fd_sc_hd__mux2_1
X_22509_ _22503_/X _22504_/X _22505_/X _22506_/X _22507_/X _22508_/X vssd1 vssd1 vccd1
+ vccd1 _22510_/A sky130_fd_sc_hd__mux4_1
XFILLER_11_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 la1_data_in[19] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14291_ _14304_/A vssd1 vssd1 vccd1 vccd1 _14302_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26277_ _20281_/X _26277_/D vssd1 vssd1 vccd1 vccd1 _26277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23489_ _27188_/Q _23495_/B vssd1 vssd1 vccd1 vccd1 _23489_/X sky130_fd_sc_hd__or2_1
XFILLER_202_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_28016_ _28016_/A _15874_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
XFILLER_7_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16030_ _16030_/A _16030_/B _16030_/C _16020_/X vssd1 vssd1 vccd1 vccd1 _16194_/C
+ sky130_fd_sc_hd__or4b_2
X_13242_ _13242_/A vssd1 vssd1 vccd1 vccd1 _27034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25228_ _25228_/A _25228_/B vssd1 vssd1 vccd1 vccd1 _25229_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25159_ _27695_/Q _25142_/X _25158_/Y _25132_/X vssd1 vssd1 vccd1 vccd1 _27695_/D
+ sky130_fd_sc_hd__o211a_1
X_13173_ _13205_/A vssd1 vssd1 vccd1 vccd1 _13199_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_151_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17981_ _17972_/X _17975_/X _17980_/X _17932_/X vssd1 vssd1 vccd1 vccd1 _17992_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19720_ _19710_/X _19711_/X _19712_/X _19713_/X _19714_/X _19715_/X vssd1 vssd1 vccd1
+ vccd1 _19721_/A sky130_fd_sc_hd__mux4_1
XFILLER_46_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16932_ _27596_/Q vssd1 vssd1 vccd1 vccd1 _18443_/A sky130_fd_sc_hd__clkinv_2
XFILLER_133_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19651_ _19651_/A vssd1 vssd1 vccd1 vccd1 _19651_/X sky130_fd_sc_hd__clkbuf_1
X_16863_ _16862_/A _16862_/B _16646_/B vssd1 vssd1 vccd1 vccd1 _16863_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18602_ _25358_/A vssd1 vssd1 vccd1 vccd1 _25625_/S sky130_fd_sc_hd__buf_2
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15814_ _13133_/X _26092_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15815_/A sky130_fd_sc_hd__mux2_1
X_19582_ _19582_/A vssd1 vssd1 vccd1 vccd1 _19582_/X sky130_fd_sc_hd__clkbuf_1
X_16794_ _16110_/A _24305_/A _16559_/A vssd1 vssd1 vccd1 vccd1 _16831_/A sky130_fd_sc_hd__o21ai_1
XFILLER_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18533_ _26839_/Q _26807_/Q _26775_/Q _26743_/Q _17832_/X _17835_/X vssd1 vssd1 vccd1
+ vccd1 _18533_/X sky130_fd_sc_hd__mux4_1
X_15745_ _15745_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15745_/Y sky130_fd_sc_hd__nor2_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _27818_/Q _12965_/B vssd1 vssd1 vccd1 vccd1 _12958_/A sky130_fd_sc_hd__and2_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18464_ _18461_/X _18463_/X _18488_/S vssd1 vssd1 vccd1 vccd1 _18464_/X sky130_fd_sc_hd__mux2_2
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15676_ _13190_/X _26146_/Q _15678_/S vssd1 vssd1 vccd1 vccd1 _15677_/A sky130_fd_sc_hd__mux2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _26818_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_282 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17415_ _27387_/Q _27386_/Q _27385_/Q _27384_/Q vssd1 vssd1 vccd1 vccd1 _17418_/A
+ sky130_fd_sc_hd__or4_1
X_14627_ _26585_/Q _14615_/X _14624_/X _14626_/Y vssd1 vssd1 vccd1 vccd1 _26585_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA_293 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18395_ _18395_/A vssd1 vssd1 vccd1 vccd1 _18488_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _17344_/X _17345_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17346_/X sky130_fd_sc_hd__mux2_2
XFILLER_147_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14558_ _15718_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14558_/Y sky130_fd_sc_hd__nor2_1
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _26954_/Q _13487_/X _13505_/X _13508_/Y vssd1 vssd1 vccd1 vccd1 _26954_/D
+ sky130_fd_sc_hd__a31o_1
X_17277_ _17338_/A vssd1 vssd1 vccd1 vccd1 _17277_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _16442_/A vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__clkbuf_2
X_27997__463 vssd1 vssd1 vccd1 vccd1 _27997__463/HI _27997_/A sky130_fd_sc_hd__conb_1
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19016_ _26689_/Q _26657_/Q _26625_/Q _26593_/Q _19015_/X _18939_/X vssd1 vssd1 vccd1
+ vccd1 _19016_/X sky130_fd_sc_hd__mux4_2
X_16228_ _26050_/Q _16235_/B _16233_/C vssd1 vssd1 vccd1 vccd1 _16228_/X sky130_fd_sc_hd__and3_1
XFILLER_161_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _16191_/B vssd1 vssd1 vccd1 vccd1 _16233_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_575 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19918_ _19988_/A vssd1 vssd1 vccd1 vccd1 _19918_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19849_ _19849_/A vssd1 vssd1 vccd1 vccd1 _19849_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_450 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22860_ _22860_/A vssd1 vssd1 vccd1 vccd1 _22860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21811_ _21827_/A vssd1 vssd1 vccd1 vccd1 _21811_/X sky130_fd_sc_hd__clkbuf_1
X_22791_ _22783_/X _22784_/X _22785_/X _22786_/X _22788_/X _22790_/X vssd1 vssd1 vccd1
+ vccd1 _22792_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_529 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24530_ _24551_/S vssd1 vssd1 vccd1 vccd1 _24545_/S sky130_fd_sc_hd__clkbuf_2
X_21742_ _22087_/A vssd1 vssd1 vccd1 vccd1 _21813_/A sky130_fd_sc_hd__buf_2
XFILLER_145_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24461_ _27628_/Q _24467_/B vssd1 vssd1 vccd1 vccd1 _24462_/A sky130_fd_sc_hd__and2_1
X_21673_ _21739_/A vssd1 vssd1 vccd1 vccd1 _21673_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23412_ _23416_/A _23416_/B _23507_/B vssd1 vssd1 vccd1 vccd1 _23413_/A sky130_fd_sc_hd__or3b_1
X_26200_ _20019_/X _26200_/D vssd1 vssd1 vccd1 vccd1 _26200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20624_ _20672_/A vssd1 vssd1 vccd1 vccd1 _20624_/X sky130_fd_sc_hd__clkbuf_2
X_27180_ _27180_/CLK _27180_/D vssd1 vssd1 vccd1 vccd1 _27180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24392_ _24392_/A _24400_/B vssd1 vssd1 vccd1 vccd1 _24393_/A sky130_fd_sc_hd__and2_1
XFILLER_132_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26131_ _19773_/X _26131_/D vssd1 vssd1 vccd1 vccd1 _26131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23343_ _27755_/Q vssd1 vssd1 vccd1 vccd1 _24733_/A sky130_fd_sc_hd__clkinv_2
X_20555_ _20587_/A vssd1 vssd1 vccd1 vccd1 _20555_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26062_ _26062_/CLK _26062_/D vssd1 vssd1 vccd1 vccd1 _26062_/Q sky130_fd_sc_hd__dfxtp_1
X_23274_ _27725_/Q _23271_/Y _23256_/Y input50/X _23273_/Y vssd1 vssd1 vccd1 vccd1
+ _23275_/D sky130_fd_sc_hd__a221o_1
X_20486_ _20480_/X _20481_/X _20482_/X _20483_/X _20484_/X _20485_/X vssd1 vssd1 vccd1
+ vccd1 _20487_/A sky130_fd_sc_hd__mux4_1
X_25013_ _25102_/S vssd1 vssd1 vccd1 vccd1 _25047_/S sky130_fd_sc_hd__clkbuf_2
X_22225_ _22213_/X _22214_/X _22215_/X _22216_/X _22217_/X _22218_/X vssd1 vssd1 vccd1
+ vccd1 _22226_/A sky130_fd_sc_hd__mux4_1
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22156_ _22156_/A vssd1 vssd1 vccd1 vccd1 _22156_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21107_ _21093_/X _21094_/X _21095_/X _21096_/X _21097_/X _21098_/X vssd1 vssd1 vccd1
+ vccd1 _21108_/A sky130_fd_sc_hd__mux4_1
XFILLER_154_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22087_ _22087_/A vssd1 vssd1 vccd1 vccd1 _22161_/A sky130_fd_sc_hd__buf_2
X_26964_ _22680_/X _26964_/D vssd1 vssd1 vccd1 vccd1 _26964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21038_ _21038_/A vssd1 vssd1 vccd1 vccd1 _21038_/X sky130_fd_sc_hd__clkbuf_1
X_25915_ _26016_/CLK _25915_/D vssd1 vssd1 vccd1 vccd1 _25915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26895_ _22442_/X _26895_/D vssd1 vssd1 vccd1 vccd1 _26895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _26840_/Q _13844_/X _13855_/X _13859_/Y vssd1 vssd1 vccd1 vccd1 _26840_/D
+ sky130_fd_sc_hd__a31o_1
X_25846_ _25878_/CLK _25846_/D vssd1 vssd1 vccd1 vccd1 _25846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25777_ _17482_/X _27844_/Q _25779_/S vssd1 vssd1 vccd1 vccd1 _25778_/A sky130_fd_sc_hd__mux2_1
X_13791_ _26864_/Q _13778_/X _13780_/X _13790_/Y vssd1 vssd1 vccd1 vccd1 _26864_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22989_ _22974_/X _22976_/X _22978_/X _22980_/X _22981_/X _22982_/X vssd1 vssd1 vccd1
+ vccd1 _22990_/A sky130_fd_sc_hd__mux4_1
X_15530_ _13184_/X _26211_/Q _15534_/S vssd1 vssd1 vccd1 vccd1 _15531_/A sky130_fd_sc_hd__mux2_1
X_27516_ _27706_/CLK _27516_/D vssd1 vssd1 vccd1 vccd1 _27516_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24728_ _27192_/Q _25474_/A vssd1 vssd1 vccd1 vccd1 _24728_/X sky130_fd_sc_hd__or2_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15461_ _15461_/A vssd1 vssd1 vccd1 vccd1 _26242_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27447_ _27447_/CLK _27447_/D vssd1 vssd1 vccd1 vccd1 _27447_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24659_ _24635_/B _24643_/X _24658_/X _24650_/X vssd1 vssd1 vccd1 vccd1 _27582_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ _25358_/B vssd1 vssd1 vccd1 vccd1 _17250_/S sky130_fd_sc_hd__clkbuf_2
X_14412_ _14412_/A _14412_/B vssd1 vssd1 vccd1 vccd1 _14412_/Y sky130_fd_sc_hd__nor2_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18180_ _18057_/X _18176_/X _18179_/X _18062_/X vssd1 vssd1 vccd1 vccd1 _18180_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27378_ _27672_/CLK _27378_/D vssd1 vssd1 vccd1 vccd1 _27378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15392_ _15392_/A vssd1 vssd1 vccd1 vccd1 _15401_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_184_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ _27836_/Q _27140_/Q _25885_/Q _25853_/Q _17081_/X _17130_/X vssd1 vssd1 vccd1
+ vccd1 _17131_/X sky130_fd_sc_hd__mux4_1
X_14343_ _26677_/Q _14337_/X _14329_/X _14342_/Y vssd1 vssd1 vccd1 vccd1 _26677_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26329_ _20463_/X _26329_/D vssd1 vssd1 vccd1 vccd1 _26329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14274_ _14361_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14274_/Y sky130_fd_sc_hd__nor2_1
X_17062_ _17385_/S vssd1 vssd1 vccd1 vccd1 _17112_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16013_ _27480_/Q _27267_/Q vssd1 vssd1 vccd1 vccd1 _16030_/B sky130_fd_sc_hd__xor2_1
X_13225_ _27273_/Q _13231_/B vssd1 vssd1 vccd1 vccd1 _13225_/X sky130_fd_sc_hd__and2_1
XFILLER_12_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13156_ _14766_/A vssd1 vssd1 vccd1 vccd1 _13156_/X sky130_fd_sc_hd__clkbuf_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_426 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _18392_/A vssd1 vssd1 vccd1 vccd1 _17964_/X sky130_fd_sc_hd__buf_2
X_13087_ _13241_/S vssd1 vssd1 vccd1 vccd1 _13112_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19703_ _19703_/A vssd1 vssd1 vccd1 vccd1 _19703_/X sky130_fd_sc_hd__clkbuf_1
X_16915_ _16915_/A _16915_/B vssd1 vssd1 vccd1 vccd1 _16915_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_66_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater406 _26047_/CLK vssd1 vssd1 vccd1 vccd1 _27312_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater417 _25958_/CLK vssd1 vssd1 vccd1 vccd1 _27333_/CLK sky130_fd_sc_hd__clkbuf_1
X_17895_ _17888_/X _17891_/X _17893_/X _17894_/X vssd1 vssd1 vccd1 vccd1 _17895_/X
+ sky130_fd_sc_hd__o211a_1
Xrepeater428 _26053_/CLK vssd1 vssd1 vccd1 vccd1 _27325_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19634_ _19634_/A vssd1 vssd1 vccd1 vccd1 _19634_/X sky130_fd_sc_hd__clkbuf_1
X_16846_ _16845_/Y _16073_/C _25908_/Q vssd1 vssd1 vccd1 vccd1 _16846_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_93_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19565_ _19563_/X _19564_/X _19565_/S vssd1 vssd1 vccd1 vccd1 _19565_/X sky130_fd_sc_hd__mux2_1
X_16777_ _16750_/X _16751_/Y _16766_/X _16844_/B vssd1 vssd1 vccd1 vccd1 _16777_/X
+ sky130_fd_sc_hd__a31o_1
X_13989_ _14361_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13989_/Y sky130_fd_sc_hd__nor2_1
X_18516_ _18516_/A _17910_/X vssd1 vssd1 vccd1 vccd1 _18516_/X sky130_fd_sc_hd__or2b_1
X_15728_ _15728_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15728_/Y sky130_fd_sc_hd__nor2_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19496_ _19496_/A vssd1 vssd1 vccd1 vccd1 _26069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18447_ _27818_/Q _26579_/Q _26451_/Q _26131_/Q _17899_/X _17997_/X vssd1 vssd1 vccd1
+ vccd1 _18447_/X sky130_fd_sc_hd__mux4_1
X_15659_ _13144_/X _26154_/Q _15667_/S vssd1 vssd1 vccd1 vccd1 _15660_/A sky130_fd_sc_hd__mux2_1
X_18378_ _18376_/X _18377_/X _18378_/S vssd1 vssd1 vccd1 vccd1 _18378_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17329_ _17277_/X _17329_/B vssd1 vssd1 vccd1 vccd1 _17329_/X sky130_fd_sc_hd__and2b_1
XFILLER_119_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20340_ _20340_/A vssd1 vssd1 vccd1 vccd1 _20413_/A sky130_fd_sc_hd__buf_2
XFILLER_88_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20271_ _20336_/A vssd1 vssd1 vccd1 vccd1 _20271_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22010_ _22010_/A vssd1 vssd1 vccd1 vccd1 _22010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_597 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23961_ _25933_/Q _25999_/Q _25832_/Q _26031_/Q _23946_/X _23929_/X vssd1 vssd1 vccd1
+ vccd1 _23961_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25700_ _25700_/A vssd1 vssd1 vccd1 vccd1 _25700_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22912_ _22944_/A vssd1 vssd1 vccd1 vccd1 _22912_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26680_ _21696_/X _26680_/D vssd1 vssd1 vccd1 vccd1 _26680_/Q sky130_fd_sc_hd__dfxtp_1
X_23892_ _27080_/Q _27112_/Q _23892_/S vssd1 vssd1 vccd1 vccd1 _23892_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22843_ _22837_/X _22838_/X _22839_/X _22840_/X _22841_/X _22842_/X vssd1 vssd1 vccd1
+ vccd1 _22844_/A sky130_fd_sc_hd__mux4_1
X_25631_ _23025_/X _23026_/X _23027_/X _23028_/X _23029_/X _23030_/X vssd1 vssd1 vccd1
+ vccd1 _25632_/A sky130_fd_sc_hd__mux4_1
XFILLER_186_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25562_ _25560_/X _25283_/B _25561_/X _25543_/X vssd1 vssd1 vccd1 vccd1 _25562_/X
+ sky130_fd_sc_hd__a211o_1
X_22774_ _22774_/A vssd1 vssd1 vccd1 vccd1 _22774_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27301_ _27789_/CLK _27301_/D vssd1 vssd1 vccd1 vccd1 _27301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21725_ _21725_/A vssd1 vssd1 vccd1 vccd1 _21725_/X sky130_fd_sc_hd__clkbuf_2
X_24513_ _27605_/Q _24554_/B vssd1 vssd1 vccd1 vccd1 _24514_/A sky130_fd_sc_hd__and2_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25493_ _25553_/A vssd1 vssd1 vccd1 vccd1 _25493_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27232_ _27232_/CLK _27232_/D vssd1 vssd1 vccd1 vccd1 _27232_/Q sky130_fd_sc_hd__dfxtp_1
X_21656_ _21656_/A vssd1 vssd1 vccd1 vccd1 _21656_/X sky130_fd_sc_hd__clkbuf_1
X_24444_ _24444_/A vssd1 vssd1 vccd1 vccd1 _27499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20607_ _20607_/A vssd1 vssd1 vccd1 vccd1 _20607_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27163_ _27574_/CLK _27163_/D vssd1 vssd1 vccd1 vccd1 _27163_/Q sky130_fd_sc_hd__dfxtp_1
X_24375_ _24375_/A vssd1 vssd1 vccd1 vccd1 _27469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21587_ _21635_/A vssd1 vssd1 vccd1 vccd1 _21587_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26114_ _19709_/X _26114_/D vssd1 vssd1 vccd1 vccd1 _26114_/Q sky130_fd_sc_hd__dfxtp_1
X_23326_ input67/X input68/X input69/X input70/X vssd1 vssd1 vccd1 vccd1 _23332_/C
+ sky130_fd_sc_hd__or4_1
X_20538_ _20586_/A vssd1 vssd1 vccd1 vccd1 _20538_/X sky130_fd_sc_hd__clkbuf_2
X_27094_ _27094_/CLK _27094_/D vssd1 vssd1 vccd1 vccd1 _27094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23257_ _27722_/Q vssd1 vssd1 vccd1 vccd1 _23257_/Y sky130_fd_sc_hd__inv_2
X_26045_ _27358_/CLK _26045_/D vssd1 vssd1 vccd1 vccd1 _26045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_520 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20469_ _20501_/A vssd1 vssd1 vccd1 vccd1 _20469_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13010_ _13010_/A vssd1 vssd1 vccd1 vccd1 _27794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22208_ _22208_/A vssd1 vssd1 vccd1 vccd1 _22208_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_669 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23188_ _23188_/A vssd1 vssd1 vccd1 vccd1 _27131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22139_ _22125_/X _22126_/X _22127_/X _22128_/X _22129_/X _22130_/X vssd1 vssd1 vccd1
+ vccd1 _22140_/A sky130_fd_sc_hd__mux4_1
XFILLER_121_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27996_ _27996_/A _15885_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_95_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26947_ _22624_/X _26947_/D vssd1 vssd1 vccd1 vccd1 _26947_/Q sky130_fd_sc_hd__dfxtp_1
X_14961_ _14975_/A vssd1 vssd1 vccd1 vccd1 _14966_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_897 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16700_ _16700_/A _16700_/B vssd1 vssd1 vccd1 vccd1 _16700_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_43_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13912_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13912_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17680_ _27409_/Q vssd1 vssd1 vccd1 vccd1 _17680_/X sky130_fd_sc_hd__clkbuf_2
X_26878_ _22382_/X _26878_/D vssd1 vssd1 vccd1 vccd1 _26878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14892_ _14718_/X _26487_/Q _14896_/S vssd1 vssd1 vccd1 vccd1 _14893_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16631_ _16631_/A _16631_/B vssd1 vssd1 vccd1 vccd1 _16631_/Y sky130_fd_sc_hd__xnor2_1
X_13843_ _26844_/Q _13832_/X _13833_/X _13842_/Y vssd1 vssd1 vccd1 vccd1 _26844_/D
+ sky130_fd_sc_hd__a31o_1
X_25829_ _27094_/CLK _25829_/D vssd1 vssd1 vccd1 vccd1 _25829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19350_ _19419_/A _19350_/B vssd1 vssd1 vccd1 vccd1 _19350_/X sky130_fd_sc_hd__or2_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16562_ _16648_/C _16570_/B vssd1 vssd1 vccd1 vccd1 _16652_/B sky130_fd_sc_hd__nor2_1
XFILLER_16_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13774_ _13868_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13774_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18301_ _18458_/A vssd1 vssd1 vccd1 vccd1 _18301_/X sky130_fd_sc_hd__buf_2
XFILLER_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15513_ _15513_/A vssd1 vssd1 vccd1 vccd1 _26219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19281_ _26156_/Q _26092_/Q _27020_/Q _26988_/Q _19165_/X _19188_/X vssd1 vssd1 vccd1
+ vccd1 _19282_/B sky130_fd_sc_hd__mux4_1
XFILLER_71_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ _16809_/B _16493_/B _16493_/C vssd1 vssd1 vccd1 vccd1 _16494_/B sky130_fd_sc_hd__and3_1
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18232_ _18162_/X _18231_/X _18211_/X vssd1 vssd1 vccd1 vccd1 _18232_/X sky130_fd_sc_hd__o21a_1
X_15444_ _15444_/A vssd1 vssd1 vccd1 vccd1 _26250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18163_ _26278_/Q _26246_/Q _26214_/Q _26182_/Q _18044_/X _18068_/X vssd1 vssd1 vccd1
+ vccd1 _18163_/X sky130_fd_sc_hd__mux4_2
X_15375_ _14766_/X _26280_/Q _15379_/S vssd1 vssd1 vccd1 vccd1 _15376_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ _27203_/Q _17113_/X _17128_/S vssd1 vssd1 vccd1 vccd1 _17115_/A sky130_fd_sc_hd__mux2_1
X_14326_ _26682_/Q _14322_/X _14248_/B _14325_/Y vssd1 vssd1 vccd1 vccd1 _26682_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18094_ _26275_/Q _26243_/Q _26211_/Q _26179_/Q _17801_/X _17805_/X vssd1 vssd1 vccd1
+ vccd1 _18094_/X sky130_fd_sc_hd__mux4_2
XFILLER_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17045_ _16998_/X _17044_/X _17033_/X vssd1 vssd1 vccd1 vccd1 _17045_/X sky130_fd_sc_hd__a21bo_1
X_14257_ _14257_/A vssd1 vssd1 vccd1 vccd1 _14311_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ _27276_/Q _13237_/B vssd1 vssd1 vccd1 vccd1 _13208_/X sky130_fd_sc_hd__and2_2
X_14188_ _26733_/Q _14186_/X _14181_/X _14187_/Y vssd1 vssd1 vccd1 vccd1 _26733_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ _14756_/A vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__buf_2
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18996_ _19431_/A vssd1 vssd1 vccd1 vccd1 _18996_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater203 _27076_/CLK vssd1 vssd1 vccd1 vccd1 _26020_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _18028_/A _17947_/B _17947_/C vssd1 vssd1 vccd1 vccd1 _17948_/A sky130_fd_sc_hd__and3_1
Xrepeater214 _27232_/CLK vssd1 vssd1 vccd1 vccd1 _27826_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater225 _26065_/CLK vssd1 vssd1 vccd1 vccd1 _27332_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater236 _27729_/CLK vssd1 vssd1 vccd1 vccd1 _27737_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater247 _27726_/CLK vssd1 vssd1 vccd1 vccd1 _27747_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater258 _27612_/CLK vssd1 vssd1 vccd1 vccd1 _27529_/CLK sky130_fd_sc_hd__clkbuf_1
X_17878_ _26395_/Q _26363_/Q _26331_/Q _26299_/Q _17877_/X _17848_/X vssd1 vssd1 vccd1
+ vccd1 _17878_/X sky130_fd_sc_hd__mux4_1
Xrepeater269 _27589_/CLK vssd1 vssd1 vccd1 vccd1 _27174_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16829_ _16648_/X _16650_/B _16565_/A vssd1 vssd1 vccd1 vccd1 _16829_/X sky130_fd_sc_hd__o21ba_1
X_19617_ _19605_/X _19606_/X _19607_/X _19608_/X _19609_/X _19610_/X vssd1 vssd1 vccd1
+ vccd1 _19618_/A sky130_fd_sc_hd__mux4_1
XFILLER_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19548_ _19542_/X _19544_/X _19547_/X _18895_/A _19469_/X vssd1 vssd1 vccd1 vccd1
+ _19549_/C sky130_fd_sc_hd__a221o_1
XFILLER_59_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19479_ _27820_/Q _26581_/Q _26453_/Q _26133_/Q _19414_/X _18831_/X vssd1 vssd1 vccd1
+ vccd1 _19479_/X sky130_fd_sc_hd__mux4_1
XFILLER_181_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21510_ _21510_/A vssd1 vssd1 vccd1 vccd1 _21510_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22490_ _22522_/A vssd1 vssd1 vccd1 vccd1 _22490_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21441_ _21427_/X _21428_/X _21429_/X _21430_/X _21431_/X _21432_/X vssd1 vssd1 vccd1
+ vccd1 _21442_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24160_ _27457_/Q _24162_/B vssd1 vssd1 vccd1 vccd1 _24161_/A sky130_fd_sc_hd__and2_1
XFILLER_175_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21372_ _21372_/A vssd1 vssd1 vccd1 vccd1 _21372_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23111_ _23167_/A vssd1 vssd1 vccd1 vccd1 _23180_/S sky130_fd_sc_hd__buf_2
XFILLER_163_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20323_ _20323_/A vssd1 vssd1 vccd1 vccd1 _20323_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24091_ _27394_/Q _24095_/B vssd1 vssd1 vccd1 vccd1 _24092_/A sky130_fd_sc_hd__and2_1
XFILLER_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23042_ _27067_/Q _17680_/X _23048_/S vssd1 vssd1 vccd1 vccd1 _23043_/A sky130_fd_sc_hd__mux2_1
X_20254_ _20340_/A vssd1 vssd1 vccd1 vccd1 _20323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27850_ _27850_/CLK _27850_/D vssd1 vssd1 vccd1 vccd1 _27850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20185_ _20250_/A vssd1 vssd1 vccd1 vccd1 _20185_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26801_ _22118_/X _26801_/D vssd1 vssd1 vccd1 vccd1 _26801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27781_ _27781_/CLK _27781_/D vssd1 vssd1 vccd1 vccd1 _27781_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24993_ _25914_/Q _25980_/Q _25813_/Q _26012_/Q _24974_/X _24983_/X vssd1 vssd1 vccd1
+ vccd1 _24993_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26732_ _21874_/X _26732_/D vssd1 vssd1 vccd1 vccd1 _26732_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23944_ _23991_/A vssd1 vssd1 vccd1 vccd1 _23944_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26663_ _21628_/X _26663_/D vssd1 vssd1 vccd1 vccd1 _26663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23875_ _25924_/Q _25990_/Q _25823_/Q _26022_/Q _23852_/X _23835_/X vssd1 vssd1 vccd1
+ vccd1 _23875_/X sky130_fd_sc_hd__mux4_1
XFILLER_189_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25614_ _24969_/A _18606_/X _25611_/Y _25613_/X _25592_/X vssd1 vssd1 vccd1 vccd1
+ _27784_/D sky130_fd_sc_hd__a221oi_1
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22826_ _22858_/A vssd1 vssd1 vccd1 vccd1 _22826_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26594_ _21388_/X _26594_/D vssd1 vssd1 vccd1 vccd1 _26594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25545_ _24780_/A _25534_/X _25541_/Y _25544_/X _25527_/X vssd1 vssd1 vccd1 vccd1
+ _27771_/D sky130_fd_sc_hd__a221oi_1
XFILLER_197_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22757_ _22751_/X _22752_/X _22753_/X _22754_/X _22755_/X _22756_/X vssd1 vssd1 vccd1
+ vccd1 _22758_/A sky130_fd_sc_hd__mux4_1
XFILLER_73_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21708_ _21740_/A vssd1 vssd1 vccd1 vccd1 _21708_/X sky130_fd_sc_hd__clkbuf_1
X_13490_ _13889_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22688_ _22688_/A vssd1 vssd1 vccd1 vccd1 _22688_/X sky130_fd_sc_hd__clkbuf_1
X_25476_ _25456_/X _25461_/X _25462_/X _24854_/B _25463_/X vssd1 vssd1 vccd1 vccd1
+ _25476_/X sky130_fd_sc_hd__o311a_1
X_27215_ _27422_/CLK _27215_/D vssd1 vssd1 vccd1 vccd1 _27215_/Q sky130_fd_sc_hd__dfxtp_1
X_21639_ _21631_/X _21632_/X _21633_/X _21634_/X _21635_/X _21636_/X vssd1 vssd1 vccd1
+ vccd1 _21640_/A sky130_fd_sc_hd__mux4_1
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24427_ _27613_/Q _24433_/B vssd1 vssd1 vccd1 vccd1 _24428_/A sky130_fd_sc_hd__and2_1
XFILLER_176_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27146_ _27844_/CLK _27146_/D vssd1 vssd1 vccd1 vccd1 _27146_/Q sky130_fd_sc_hd__dfxtp_1
X_15160_ _26375_/Q _13379_/X _15162_/S vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24358_ _24358_/A vssd1 vssd1 vccd1 vccd1 _27461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14111_ _26761_/Q _14104_/X _14107_/X _14110_/Y vssd1 vssd1 vccd1 vccd1 _26761_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_181_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23309_ _23309_/A _23309_/B _23309_/C vssd1 vssd1 vccd1 vccd1 _23321_/C sky130_fd_sc_hd__or3_1
X_15091_ _15091_/A vssd1 vssd1 vccd1 vccd1 _26406_/D sky130_fd_sc_hd__clkbuf_1
X_27077_ _27077_/CLK _27077_/D vssd1 vssd1 vccd1 vccd1 _27077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24289_ _24330_/A vssd1 vssd1 vccd1 vccd1 _24317_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14042_ _14090_/A vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26028_ _27095_/CLK _26028_/D vssd1 vssd1 vccd1 vccd1 _26028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ _26939_/Q _26907_/Q _26875_/Q _26843_/Q _18788_/X _18790_/X vssd1 vssd1 vccd1
+ vccd1 _18850_/X sky130_fd_sc_hd__mux4_2
XFILLER_192_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17801_ _18085_/A vssd1 vssd1 vccd1 vccd1 _17801_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18781_ _18923_/A vssd1 vssd1 vccd1 vccd1 _19227_/A sky130_fd_sc_hd__buf_2
X_27979_ _27979_/A _15905_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_15993_ _16034_/A vssd1 vssd1 vccd1 vccd1 _16242_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17732_ _25929_/Q _17731_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17733_/A sky130_fd_sc_hd__mux2_1
X_14944_ _14944_/A vssd1 vssd1 vccd1 vccd1 _26464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17663_ _17511_/X _25902_/Q _17667_/S vssd1 vssd1 vccd1 vccd1 _17664_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_473 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14875_ _26494_/Q _13408_/X _14879_/S vssd1 vssd1 vccd1 vccd1 _14876_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19402_ _26545_/Q _26513_/Q _26481_/Q _27057_/Q _19401_/X _19287_/X vssd1 vssd1 vccd1
+ vccd1 _19402_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16614_ _16616_/A _16616_/B vssd1 vssd1 vccd1 vccd1 _16614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _26851_/Q _13819_/X _13820_/X _13825_/Y vssd1 vssd1 vccd1 vccd1 _26851_/D
+ sky130_fd_sc_hd__a31o_1
X_17594_ _17594_/A vssd1 vssd1 vccd1 vccd1 _25871_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19333_ _26542_/Q _26510_/Q _26478_/Q _27054_/Q _19242_/X _19287_/X vssd1 vssd1 vccd1
+ vccd1 _19333_/X sky130_fd_sc_hd__mux4_1
X_16545_ _16815_/B _16545_/B vssd1 vssd1 vccd1 vccd1 _16545_/X sky130_fd_sc_hd__and2_1
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _13938_/A _13759_/B vssd1 vssd1 vccd1 vccd1 _13757_/Y sky130_fd_sc_hd__nor2_1
X_19264_ _26411_/Q _26379_/Q _26347_/Q _26315_/Q _19170_/X _19240_/X vssd1 vssd1 vccd1
+ vccd1 _19264_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16476_ _16786_/B _16476_/B vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__nand2_1
X_13688_ _26902_/Q _13682_/X _13676_/X _13687_/Y vssd1 vssd1 vccd1 vccd1 _26902_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_188_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18215_ _26408_/Q _26376_/Q _26344_/Q _26312_/Q _18189_/X _18214_/X vssd1 vssd1 vccd1
+ vccd1 _18215_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15427_ _26257_/Q _13347_/X _15429_/S vssd1 vssd1 vccd1 vccd1 _15428_/A sky130_fd_sc_hd__mux2_1
X_19195_ _19191_/X _19193_/X _19194_/X vssd1 vssd1 vccd1 vccd1 _19195_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_431 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_28022__488 vssd1 vssd1 vccd1 vccd1 _28022__488/HI _28022_/A sky130_fd_sc_hd__conb_1
XFILLER_157_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18146_ _18146_/A _18146_/B _18146_/C vssd1 vssd1 vccd1 vccd1 _18147_/A sky130_fd_sc_hd__and3_1
XFILLER_191_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ _15358_/A vssd1 vssd1 vccd1 vccd1 _26288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ _14548_/A vssd1 vssd1 vccd1 vccd1 _14365_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18077_ _18146_/A _18077_/B _18077_/C vssd1 vssd1 vccd1 vccd1 _18078_/A sky130_fd_sc_hd__and3_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15289_ _26318_/Q _13357_/X _15295_/S vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17028_ _27828_/Q _27132_/Q _25877_/Q _25845_/Q _17015_/X _16989_/X vssd1 vssd1 vccd1
+ vccd1 _17028_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _19004_/A _18979_/B vssd1 vssd1 vccd1 vccd1 _18979_/X sky130_fd_sc_hd__or2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21990_ _21990_/A vssd1 vssd1 vccd1 vccd1 _21990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20941_ _20941_/A vssd1 vssd1 vccd1 vccd1 _20941_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23660_ _23660_/A vssd1 vssd1 vccd1 vccd1 _27236_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20872_ _22616_/A vssd1 vssd1 vccd1 vccd1 _21217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_476 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22611_ _22611_/A vssd1 vssd1 vccd1 vccd1 _22611_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23591_ _27776_/Q _27218_/Q _23595_/S vssd1 vssd1 vccd1 vccd1 _23592_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22542_ _22610_/A vssd1 vssd1 vccd1 vccd1 _22542_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25330_ _27514_/Q _27513_/Q _25332_/A vssd1 vssd1 vccd1 vccd1 _25330_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_201_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22473_ _22521_/A vssd1 vssd1 vccd1 vccd1 _22473_/X sky130_fd_sc_hd__clkbuf_1
X_25261_ _25261_/A _25261_/B vssd1 vssd1 vccd1 vccd1 _25261_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27000_ _22812_/X _27000_/D vssd1 vssd1 vccd1 vccd1 _27000_/Q sky130_fd_sc_hd__dfxtp_1
X_21424_ _21424_/A vssd1 vssd1 vccd1 vccd1 _21424_/X sky130_fd_sc_hd__clkbuf_1
X_24212_ _24380_/B vssd1 vssd1 vccd1 vccd1 _24233_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25192_ _25221_/A _25192_/B vssd1 vssd1 vccd1 vccd1 _25192_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24143_ _27449_/Q _24151_/B vssd1 vssd1 vccd1 vccd1 _24144_/A sky130_fd_sc_hd__and2_1
X_21355_ _21341_/X _21342_/X _21343_/X _21344_/X _21345_/X _21346_/X vssd1 vssd1 vccd1
+ vccd1 _21356_/A sky130_fd_sc_hd__mux4_1
XFILLER_190_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20306_ _20322_/A vssd1 vssd1 vccd1 vccd1 _20306_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24074_ _24186_/A vssd1 vssd1 vccd1 vccd1 _24119_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_190_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21286_ _21302_/A vssd1 vssd1 vccd1 vccd1 _21286_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23025_ _25635_/A vssd1 vssd1 vccd1 vccd1 _23025_/X sky130_fd_sc_hd__clkbuf_1
X_20237_ _20237_/A vssd1 vssd1 vccd1 vccd1 _20237_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27833_ _27833_/CLK _27833_/D vssd1 vssd1 vccd1 vccd1 _27833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20168_ _20340_/A vssd1 vssd1 vccd1 vccd1 _20237_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27764_ _27772_/CLK _27764_/D vssd1 vssd1 vccd1 vccd1 _27764_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24976_ _25912_/Q _25978_/Q _25811_/Q _26010_/Q _24974_/X _24975_/X vssd1 vssd1 vccd1
+ vccd1 _24976_/X sky130_fd_sc_hd__mux4_1
X_12990_ _27803_/Q _12998_/B vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__and2_1
XFILLER_58_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20099_ _20164_/A vssd1 vssd1 vccd1 vccd1 _20099_/X sky130_fd_sc_hd__clkbuf_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26715_ _21816_/X _26715_/D vssd1 vssd1 vccd1 vccd1 _26715_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23927_ _23896_/X _23925_/X _23926_/X _23911_/X vssd1 vssd1 vccd1 vccd1 _27288_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27695_ _27695_/CLK _27695_/D vssd1 vssd1 vccd1 vccd1 _27695_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26646_ _21572_/X _26646_/D vssd1 vssd1 vccd1 vccd1 _26646_/Q sky130_fd_sc_hd__dfxtp_1
X_14660_ _26573_/Q _14658_/X _14653_/X _14659_/Y vssd1 vssd1 vccd1 vccd1 _26573_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23858_ _24047_/S vssd1 vssd1 vccd1 vccd1 _23893_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13882_/A _13621_/B vssd1 vssd1 vccd1 vccd1 _13611_/Y sky130_fd_sc_hd__nor2_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22809_ _22857_/A vssd1 vssd1 vccd1 vccd1 _22809_/X sky130_fd_sc_hd__clkbuf_2
X_14591_ _26598_/Q _14589_/X _14579_/X _14590_/Y vssd1 vssd1 vccd1 vccd1 _26598_/D
+ sky130_fd_sc_hd__a31o_1
X_26577_ _21336_/X _26577_/D vssd1 vssd1 vccd1 vccd1 _26577_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23789_ _27069_/Q _27101_/Q _23796_/S vssd1 vssd1 vccd1 vccd1 _23789_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16330_ _16360_/A _16755_/A _16336_/B vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__a21o_1
XFILLER_197_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13542_ _13917_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25528_ _24772_/A _25504_/X _25521_/Y _25526_/X _25527_/X vssd1 vssd1 vccd1 vccd1
+ _27768_/D sky130_fd_sc_hd__a221oi_1
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16261_ _27538_/Q _16109_/A vssd1 vssd1 vccd1 vccd1 _16261_/X sky130_fd_sc_hd__or2b_1
XFILLER_158_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13473_ _27358_/Q _13063_/A _13082_/X _27326_/Q _13103_/X vssd1 vssd1 vccd1 vccd1
+ _14448_/A sky130_fd_sc_hd__a221oi_4
XFILLER_13_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25459_ _24740_/A _25431_/X _25455_/Y _25458_/X _25446_/X vssd1 vssd1 vccd1 vccd1
+ _27757_/D sky130_fd_sc_hd__a221oi_1
X_18000_ _18000_/A vssd1 vssd1 vccd1 vccd1 _18000_/X sky130_fd_sc_hd__buf_2
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15212_ _14740_/X _26352_/Q _15212_/S vssd1 vssd1 vccd1 vccd1 _15213_/A sky130_fd_sc_hd__mux2_1
XFILLER_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16192_ _27521_/Q _15991_/A vssd1 vssd1 vccd1 vccd1 _16192_/X sky130_fd_sc_hd__or2b_1
XFILLER_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27129_ _27129_/CLK _27129_/D vssd1 vssd1 vccd1 vccd1 _27129_/Q sky130_fd_sc_hd__dfxtp_1
X_15143_ _26383_/Q _13353_/X _15151_/S vssd1 vssd1 vccd1 vccd1 _15144_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19951_ _19951_/A vssd1 vssd1 vccd1 vccd1 _19951_/X sky130_fd_sc_hd__clkbuf_1
X_15074_ _15074_/A vssd1 vssd1 vccd1 vccd1 _26414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14025_ _14497_/A vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__buf_2
X_18902_ _27796_/Q _26557_/Q _26429_/Q _26109_/Q _18900_/X _18901_/X vssd1 vssd1 vccd1
+ vccd1 _18902_/X sky130_fd_sc_hd__mux4_2
XFILLER_141_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19882_ _19898_/A vssd1 vssd1 vccd1 vccd1 _19882_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18833_ _18945_/A vssd1 vssd1 vccd1 vccd1 _19391_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18764_ _19428_/A vssd1 vssd1 vccd1 vccd1 _18969_/A sky130_fd_sc_hd__clkbuf_1
X_15976_ _15979_/A vssd1 vssd1 vccd1 vccd1 _15976_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17715_ _27420_/Q vssd1 vssd1 vccd1 vccd1 _17715_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ _14769_/X _26471_/Q _14929_/S vssd1 vssd1 vccd1 vccd1 _14928_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18695_ _18695_/A vssd1 vssd1 vccd1 vccd1 _26010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17646_ _17646_/A vssd1 vssd1 vccd1 vccd1 _25894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14858_ _14858_/A vssd1 vssd1 vccd1 vccd1 _26502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ _26858_/Q _13806_/X _13807_/X _13808_/Y vssd1 vssd1 vccd1 vccd1 _26858_/D
+ sky130_fd_sc_hd__a31o_1
X_17577_ _17577_/A vssd1 vssd1 vccd1 vccd1 _25863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14789_ _14788_/X _26529_/Q _14789_/S vssd1 vssd1 vccd1 vccd1 _14790_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19316_ _19409_/A _19316_/B vssd1 vssd1 vccd1 vccd1 _19316_/X sky130_fd_sc_hd__or2_1
XFILLER_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16528_ _25965_/Q vssd1 vssd1 vccd1 vccd1 _16528_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19247_ _19247_/A vssd1 vssd1 vccd1 vccd1 _26058_/D sky130_fd_sc_hd__clkbuf_1
X_16459_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16778_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19178_ _19250_/A _19178_/B vssd1 vssd1 vccd1 vccd1 _19178_/X sky130_fd_sc_hd__or2_1
XFILLER_118_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18129_ _18427_/A vssd1 vssd1 vccd1 vccd1 _18129_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21140_ _21140_/A vssd1 vssd1 vccd1 vccd1 _21140_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21071_ _21058_/X _21060_/X _21062_/X _21064_/X _21065_/X _21066_/X vssd1 vssd1 vccd1
+ vccd1 _21072_/A sky130_fd_sc_hd__mux4_1
X_20022_ _20009_/X _20011_/X _20013_/X _20015_/X _20016_/X _20017_/X vssd1 vssd1 vccd1
+ vccd1 _20023_/A sky130_fd_sc_hd__mux4_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24830_ _24940_/A vssd1 vssd1 vccd1 vccd1 _24838_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24761_ _27618_/Q _24758_/X _24759_/Y _24760_/X vssd1 vssd1 vccd1 vccd1 _27618_/D
+ sky130_fd_sc_hd__o211a_1
X_21973_ _21965_/X _21966_/X _21967_/X _21968_/X _21969_/X _21970_/X vssd1 vssd1 vccd1
+ vccd1 _21974_/A sky130_fd_sc_hd__mux4_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26500_ _21068_/X _26500_/D vssd1 vssd1 vccd1 vccd1 _26500_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23712_ _24954_/B _27260_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23713_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20924_ _20956_/A vssd1 vssd1 vccd1 vccd1 _20924_/X sky130_fd_sc_hd__clkbuf_1
X_27480_ _27480_/CLK _27480_/D vssd1 vssd1 vccd1 vccd1 _27480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24692_ _27178_/Q _24698_/B vssd1 vssd1 vccd1 vccd1 _24692_/X sky130_fd_sc_hd__or2_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_26431_ _20825_/X _26431_/D vssd1 vssd1 vccd1 vccd1 _26431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20855_/A vssd1 vssd1 vccd1 vccd1 _20855_/X sky130_fd_sc_hd__clkbuf_1
X_23643_ _25003_/S vssd1 vssd1 vccd1 vccd1 _23643_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26362_ _20577_/X _26362_/D vssd1 vssd1 vccd1 vccd1 _26362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23574_ _23577_/A _23574_/B vssd1 vssd1 vccd1 vccd1 _23575_/A sky130_fd_sc_hd__and2_1
X_20786_ _20770_/X _20771_/X _20772_/X _20773_/X _20775_/X _20777_/X vssd1 vssd1 vccd1
+ vccd1 _20787_/A sky130_fd_sc_hd__mux4_1
X_25313_ _25344_/A _25313_/B vssd1 vssd1 vccd1 vccd1 _25313_/Y sky130_fd_sc_hd__nand2_1
X_22525_ _22525_/A vssd1 vssd1 vccd1 vccd1 _22598_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_195_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26293_ _20331_/X _26293_/D vssd1 vssd1 vccd1 vccd1 _26293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25244_ _25266_/A _25244_/B vssd1 vssd1 vccd1 vccd1 _25245_/B sky130_fd_sc_hd__xnor2_1
X_22456_ _22521_/A vssd1 vssd1 vccd1 vccd1 _22456_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21407_ _21579_/A vssd1 vssd1 vccd1 vccd1 _21475_/A sky130_fd_sc_hd__clkbuf_2
X_22387_ _22435_/A vssd1 vssd1 vccd1 vccd1 _22387_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25175_ _25297_/A vssd1 vssd1 vccd1 vccd1 _25175_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_445 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21338_ _21338_/A vssd1 vssd1 vccd1 vccd1 _21338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24126_ _27442_/Q _24128_/B vssd1 vssd1 vccd1 vccd1 _24127_/A sky130_fd_sc_hd__and2_1
XFILLER_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21269_ _21301_/A vssd1 vssd1 vccd1 vccd1 _21269_/X sky130_fd_sc_hd__clkbuf_1
X_24057_ _27379_/Q _24061_/B vssd1 vssd1 vccd1 vccd1 _24058_/A sky130_fd_sc_hd__and2_1
XFILLER_151_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23008_ _23008_/A vssd1 vssd1 vccd1 vccd1 _23008_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27816_ _25704_/X _27816_/D vssd1 vssd1 vccd1 vccd1 _27816_/Q sky130_fd_sc_hd__dfxtp_1
X_15830_ _13172_/X _26085_/Q _15838_/S vssd1 vssd1 vccd1 vccd1 _15831_/A sky130_fd_sc_hd__mux2_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _15761_/A vssd1 vssd1 vccd1 vccd1 _15771_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_27747_ _27747_/CLK _27747_/D vssd1 vssd1 vccd1 vccd1 _27747_/Q sky130_fd_sc_hd__dfxtp_1
X_12973_ _12973_/A vssd1 vssd1 vccd1 vccd1 _27811_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24959_ _24960_/A _24960_/B vssd1 vssd1 vccd1 vccd1 _24965_/B sky130_fd_sc_hd__and2_1
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17500_ _17500_/A vssd1 vssd1 vccd1 vccd1 _25834_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14811_/S vssd1 vssd1 vccd1 vccd1 _14725_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18480_ _18480_/A _18479_/X vssd1 vssd1 vccd1 vccd1 _18480_/X sky130_fd_sc_hd__or2b_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27678_ _27678_/CLK _27678_/D vssd1 vssd1 vccd1 vccd1 _27969_/A sky130_fd_sc_hd__dfxtp_1
X_15692_ _15692_/A vssd1 vssd1 vccd1 vccd1 _26139_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17431_ _27410_/Q vssd1 vssd1 vccd1 vccd1 _17431_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26629_ _21512_/X _26629_/D vssd1 vssd1 vccd1 vccd1 _26629_/Q sky130_fd_sc_hd__dfxtp_1
X_14643_ _15716_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17362_ _25840_/Q _26039_/Q _17382_/S vssd1 vssd1 vccd1 vccd1 _17362_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14574_ _15736_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14574_/Y sky130_fd_sc_hd__nor2_1
XFILLER_202_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19101_ _26404_/Q _26372_/Q _26340_/Q _26308_/Q _19054_/X _19100_/X vssd1 vssd1 vccd1
+ vccd1 _19101_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16313_ _16353_/A _16313_/B _16313_/C vssd1 vssd1 vccd1 vccd1 _16384_/A sky130_fd_sc_hd__and3_1
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _16442_/A vssd1 vssd1 vccd1 vccd1 _13910_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_158_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17293_ _17242_/X _17292_/X _17281_/X vssd1 vssd1 vccd1 vccd1 _17293_/X sky130_fd_sc_hd__a21bo_1
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19032_ _19287_/A vssd1 vssd1 vccd1 vccd1 _19032_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16244_ _27389_/Q _16244_/B _16244_/C vssd1 vssd1 vccd1 vccd1 _16244_/X sky130_fd_sc_hd__and3_1
XFILLER_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13456_ _13456_/A vssd1 vssd1 vccd1 vccd1 _13553_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16175_ _16201_/A vssd1 vssd1 vccd1 vccd1 _16224_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_13387_ _26981_/Q _13385_/X _13399_/S vssd1 vssd1 vccd1 vccd1 _13388_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15126_ _15126_/A vssd1 vssd1 vccd1 vccd1 _26391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19934_ _19918_/X _19921_/X _19924_/X _19927_/X _19928_/X _19929_/X vssd1 vssd1 vccd1
+ vccd1 _19935_/A sky130_fd_sc_hd__mux4_1
X_15057_ _14724_/X _26421_/Q _15057_/S vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14008_ _26793_/Q _14005_/X _14001_/X _14007_/Y vssd1 vssd1 vccd1 vccd1 _26793_/D
+ sky130_fd_sc_hd__a31o_1
X_19865_ _19865_/A vssd1 vssd1 vccd1 vccd1 _19865_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18816_ _19317_/A vssd1 vssd1 vccd1 vccd1 _18816_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_505 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19796_ _19812_/A vssd1 vssd1 vccd1 vccd1 _19796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18747_ _18747_/A vssd1 vssd1 vccd1 vccd1 _26034_/D sky130_fd_sc_hd__clkbuf_1
X_15959_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15959_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18678_ _18678_/A vssd1 vssd1 vccd1 vccd1 _26003_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17629_ _17629_/A vssd1 vssd1 vccd1 vccd1 _25886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20640_ _20672_/A vssd1 vssd1 vccd1 vccd1 _20640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20571_ _20587_/A vssd1 vssd1 vccd1 vccd1 _20571_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22310_ _22310_/A vssd1 vssd1 vccd1 vccd1 _22310_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23290_ input66/X vssd1 vssd1 vccd1 vccd1 _23290_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22241_ _22229_/X _22230_/X _22231_/X _22232_/X _22233_/X _22234_/X vssd1 vssd1 vccd1
+ vccd1 _22242_/A sky130_fd_sc_hd__mux4_1
XFILLER_11_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22172_ _22172_/A vssd1 vssd1 vccd1 vccd1 _22172_/X sky130_fd_sc_hd__clkbuf_1
X_21123_ _21109_/X _21110_/X _21111_/X _21112_/X _21113_/X _21114_/X vssd1 vssd1 vccd1
+ vccd1 _21124_/A sky130_fd_sc_hd__mux4_1
X_26980_ _22742_/X _26980_/D vssd1 vssd1 vccd1 vccd1 _26980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25931_ _27126_/CLK _25931_/D vssd1 vssd1 vccd1 vccd1 _25931_/Q sky130_fd_sc_hd__dfxtp_1
X_21054_ _21054_/A vssd1 vssd1 vccd1 vccd1 _21054_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20005_ _20005_/A vssd1 vssd1 vccd1 vccd1 _20005_/X sky130_fd_sc_hd__clkbuf_1
X_25862_ _27149_/CLK _25862_/D vssd1 vssd1 vccd1 vccd1 _25862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27601_ _27601_/CLK _27601_/D vssd1 vssd1 vccd1 vccd1 _27601_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24813_ _24861_/A vssd1 vssd1 vccd1 vccd1 _24813_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_1157 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25793_ _17504_/X _27851_/Q _25801_/S vssd1 vssd1 vccd1 vccd1 _25794_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27532_ _27610_/CLK _27532_/D vssd1 vssd1 vccd1 vccd1 _27532_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24744_ _24744_/A _24970_/A vssd1 vssd1 vccd1 vccd1 _24744_/Y sky130_fd_sc_hd__nand2_1
X_21956_ _21956_/A vssd1 vssd1 vccd1 vccd1 _21956_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20955_/A vssd1 vssd1 vccd1 vccd1 _20907_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27463_ _27563_/CLK _27463_/D vssd1 vssd1 vccd1 vccd1 _27463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24675_ _27172_/Q _24685_/B vssd1 vssd1 vccd1 vccd1 _24675_/X sky130_fd_sc_hd__or2_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21887_ _21879_/X _21880_/X _21881_/X _21882_/X _21883_/X _21884_/X vssd1 vssd1 vccd1
+ vccd1 _21888_/A sky130_fd_sc_hd__mux4_1
XFILLER_43_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26414_ _20753_/X _26414_/D vssd1 vssd1 vccd1 vccd1 _26414_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23626_ _27227_/Q _25430_/B vssd1 vssd1 vccd1 vccd1 _27227_/D sky130_fd_sc_hd__nor2_1
XFILLER_14_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _20832_/X _20833_/X _20834_/X _20835_/X _20836_/X _20837_/X vssd1 vssd1 vccd1
+ vccd1 _20839_/A sky130_fd_sc_hd__mux4_1
X_27394_ _27394_/CLK _27394_/D vssd1 vssd1 vccd1 vccd1 _27394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26345_ _20521_/X _26345_/D vssd1 vssd1 vccd1 vccd1 _26345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23557_ _23560_/A _23557_/B vssd1 vssd1 vccd1 vccd1 _23558_/A sky130_fd_sc_hd__and2_1
X_20769_ _20769_/A vssd1 vssd1 vccd1 vccd1 _20769_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13310_/A vssd1 vssd1 vccd1 vccd1 _27006_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22508_ _22508_/A vssd1 vssd1 vccd1 vccd1 _22508_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _26696_/Q _14283_/X _14284_/X _14289_/Y vssd1 vssd1 vccd1 vccd1 _26696_/D
+ sky130_fd_sc_hd__a31o_1
X_26276_ _20279_/X _26276_/D vssd1 vssd1 vccd1 vccd1 _26276_/Q sky130_fd_sc_hd__dfxtp_1
X_23488_ input26/X _23482_/X _23486_/X _23487_/X vssd1 vssd1 vccd1 vccd1 _27187_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1117 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_28015_ _28015_/A _15862_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
XFILLER_183_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25227_ _27534_/Q _27502_/Q vssd1 vssd1 vccd1 vccd1 _25228_/B sky130_fd_sc_hd__or2_1
X_13241_ _27034_/Q _13240_/X _13241_/S vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__mux2_1
X_22439_ _22525_/A vssd1 vssd1 vccd1 vccd1 _22508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25158_ _25182_/A _25158_/B vssd1 vssd1 vccd1 vccd1 _25158_/Y sky130_fd_sc_hd__nand2_1
X_13172_ _14775_/A vssd1 vssd1 vccd1 vccd1 _13172_/X sky130_fd_sc_hd__buf_2
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24109_ _27402_/Q _24117_/B vssd1 vssd1 vccd1 vccd1 _24110_/A sky130_fd_sc_hd__and2_1
X_17980_ _17888_/X _17976_/X _17979_/X _17894_/X vssd1 vssd1 vccd1 vccd1 _17980_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25089_ _25087_/X _25088_/X _25103_/S vssd1 vssd1 vccd1 vccd1 _25089_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16931_ _27488_/Q vssd1 vssd1 vccd1 vccd1 _24210_/A sky130_fd_sc_hd__inv_2
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16862_ _16862_/A _16862_/B vssd1 vssd1 vccd1 vccd1 _16862_/Y sky130_fd_sc_hd__nor2_1
X_19650_ _19637_/X _19638_/X _19639_/X _19640_/X _19644_/X _19647_/X vssd1 vssd1 vccd1
+ vccd1 _19651_/A sky130_fd_sc_hd__mux4_1
X_18601_ _18601_/A vssd1 vssd1 vccd1 vccd1 _25110_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_15813_ _15813_/A vssd1 vssd1 vccd1 vccd1 _26093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19581_ _19570_/X _19572_/X _19574_/X _19576_/X _19577_/X _19578_/X vssd1 vssd1 vccd1
+ vccd1 _19582_/A sky130_fd_sc_hd__mux4_1
X_16793_ _16793_/A _16838_/A _16793_/C _16793_/D vssd1 vssd1 vccd1 vccd1 _16800_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18532_ _18530_/X _18531_/X _18532_/S vssd1 vssd1 vccd1 vccd1 _18532_/X sky130_fd_sc_hd__mux2_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _26121_/Q _15734_/X _15740_/X _15743_/Y vssd1 vssd1 vccd1 vccd1 _26121_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12956_ _13000_/A vssd1 vssd1 vccd1 vccd1 _12965_/B sky130_fd_sc_hd__clkbuf_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _26419_/Q _26387_/Q _26355_/Q _26323_/Q _18462_/X _18329_/X vssd1 vssd1 vccd1
+ vccd1 _18463_/X sky130_fd_sc_hd__mux4_1
X_15675_ _15675_/A vssd1 vssd1 vccd1 vccd1 _26147_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 _27773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_261 _26819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _27391_/Q _27390_/Q _27389_/Q _27388_/Q vssd1 vssd1 vccd1 vccd1 _17419_/B
+ sky130_fd_sc_hd__or4_1
X_14626_ _15699_/A _14631_/B vssd1 vssd1 vccd1 vccd1 _14626_/Y sky130_fd_sc_hd__nor2_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18394_ _26416_/Q _26384_/Q _26352_/Q _26320_/Q _18305_/X _18329_/X vssd1 vssd1 vccd1
+ vccd1 _18394_/X sky130_fd_sc_hd__mux4_1
XANTENNA_294 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17345_ _27093_/Q _27125_/Q _17355_/S vssd1 vssd1 vccd1 vccd1 _17345_/X sky130_fd_sc_hd__mux2_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _26611_/Q _14549_/X _14553_/X _14556_/Y vssd1 vssd1 vccd1 vccd1 _26611_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13508_ _13900_/A _13517_/B vssd1 vssd1 vccd1 vccd1 _13508_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17276_ _27848_/Q _27152_/Q _25897_/Q _25865_/Q _17264_/X _17252_/X vssd1 vssd1 vccd1
+ vccd1 _17276_/X sky130_fd_sc_hd__mux4_1
XFILLER_159_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _26631_/Q _14478_/X _14474_/X _14487_/Y vssd1 vssd1 vccd1 vccd1 _26631_/D
+ sky130_fd_sc_hd__a31o_1
X_19015_ _19317_/A vssd1 vssd1 vccd1 vccd1 _19015_/X sky130_fd_sc_hd__buf_2
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16227_ _16378_/A _16388_/A _16357_/A _16745_/A vssd1 vssd1 vccd1 vccd1 _16407_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_174_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13439_ _26968_/Q _13435_/X _13429_/X _13438_/Y vssd1 vssd1 vccd1 vccd1 _26968_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16158_ _27387_/Q vssd1 vssd1 vccd1 vccd1 _16420_/A sky130_fd_sc_hd__inv_2
XFILLER_170_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ _15109_/A vssd1 vssd1 vccd1 vccd1 _26398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16089_ _25910_/Q vssd1 vssd1 vccd1 vccd1 _16639_/A sky130_fd_sc_hd__buf_2
XFILLER_69_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19917_ _20266_/A vssd1 vssd1 vccd1 vccd1 _19988_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19848_ _19831_/X _19833_/X _19835_/X _19837_/X _19838_/X _19839_/X vssd1 vssd1 vccd1
+ vccd1 _19849_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _19779_/A vssd1 vssd1 vccd1 vccd1 _19779_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21810_ _21826_/A vssd1 vssd1 vccd1 vccd1 _21810_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22790_ _22858_/A vssd1 vssd1 vccd1 vccd1 _22790_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21741_ _22613_/A vssd1 vssd1 vccd1 vccd1 _22087_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24460_ _24460_/A vssd1 vssd1 vccd1 vccd1 _27506_/D sky130_fd_sc_hd__clkbuf_1
X_21672_ _22019_/A vssd1 vssd1 vccd1 vccd1 _21739_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23411_ _27782_/Q _23333_/Y _13244_/B _23337_/X _23410_/Y vssd1 vssd1 vccd1 vccd1
+ _23507_/B sky130_fd_sc_hd__o2111a_2
X_20623_ _20687_/A vssd1 vssd1 vccd1 vccd1 _20623_/X sky130_fd_sc_hd__clkbuf_1
X_24391_ _24538_/A vssd1 vssd1 vccd1 vccd1 _24400_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26130_ _19771_/X _26130_/D vssd1 vssd1 vccd1 vccd1 _26130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20554_ _20586_/A vssd1 vssd1 vccd1 vccd1 _20554_/X sky130_fd_sc_hd__clkbuf_2
X_23342_ _24776_/A _27249_/Q _27247_/Q _24769_/A vssd1 vssd1 vccd1 vccd1 _23361_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26061_ _27326_/CLK _26061_/D vssd1 vssd1 vccd1 vccd1 _26061_/Q sky130_fd_sc_hd__dfxtp_1
X_23273_ _23260_/Y input71/X _23272_/Y input44/X vssd1 vssd1 vccd1 vccd1 _23273_/Y
+ sky130_fd_sc_hd__o22ai_1
X_20485_ _20501_/A vssd1 vssd1 vccd1 vccd1 _20485_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25012_ _25008_/X _25010_/X _25046_/S vssd1 vssd1 vccd1 vccd1 _25012_/X sky130_fd_sc_hd__mux2_1
X_22224_ _22224_/A vssd1 vssd1 vccd1 vccd1 _22224_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22155_ _22141_/X _22142_/X _22143_/X _22144_/X _22145_/X _22146_/X vssd1 vssd1 vccd1
+ vccd1 _22156_/A sky130_fd_sc_hd__mux4_1
XFILLER_117_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21106_ _21106_/A vssd1 vssd1 vccd1 vccd1 _21106_/X sky130_fd_sc_hd__clkbuf_1
X_22086_ _22086_/A vssd1 vssd1 vccd1 vccd1 _22086_/X sky130_fd_sc_hd__clkbuf_1
X_26963_ _22678_/X _26963_/D vssd1 vssd1 vccd1 vccd1 _26963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21037_ _21023_/X _21024_/X _21025_/X _21026_/X _21027_/X _21028_/X vssd1 vssd1 vccd1
+ vccd1 _21038_/A sky130_fd_sc_hd__mux4_1
XFILLER_102_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25914_ _25980_/CLK _25914_/D vssd1 vssd1 vccd1 vccd1 _25914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26894_ _22432_/X _26894_/D vssd1 vssd1 vccd1 vccd1 _26894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_538 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25845_ _27132_/CLK _25845_/D vssd1 vssd1 vccd1 vccd1 _25845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25776_ _25776_/A vssd1 vssd1 vccd1 vccd1 _27843_/D sky130_fd_sc_hd__clkbuf_1
X_13790_ _13884_/A _13799_/B vssd1 vssd1 vccd1 vccd1 _13790_/Y sky130_fd_sc_hd__nor2_1
X_22988_ _22988_/A vssd1 vssd1 vccd1 vccd1 _22988_/X sky130_fd_sc_hd__clkbuf_1
X_27515_ _27515_/CLK _27515_/D vssd1 vssd1 vccd1 vccd1 _27515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24727_ _24771_/A vssd1 vssd1 vccd1 vccd1 _24727_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_21939_ _21930_/X _21932_/X _21934_/X _21936_/X _21937_/X _21938_/X vssd1 vssd1 vccd1
+ vccd1 _21940_/A sky130_fd_sc_hd__mux4_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15460_ _26242_/Q _13395_/X _15462_/S vssd1 vssd1 vccd1 vccd1 _15461_/A sky130_fd_sc_hd__mux2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27446_ _27568_/CLK _27446_/D vssd1 vssd1 vccd1 vccd1 _27446_/Q sky130_fd_sc_hd__dfxtp_1
X_24658_ _27166_/Q _24658_/B vssd1 vssd1 vccd1 vccd1 _24658_/X sky130_fd_sc_hd__or2_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _26651_/Q _14405_/X _14335_/B _14410_/Y vssd1 vssd1 vccd1 vccd1 _26651_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23609_ _23617_/A _23609_/B vssd1 vssd1 vccd1 vccd1 _23610_/A sky130_fd_sc_hd__and2_1
X_15391_ _15391_/A vssd1 vssd1 vccd1 vccd1 _26273_/D sky130_fd_sc_hd__clkbuf_1
X_27377_ _27377_/CLK _27377_/D vssd1 vssd1 vccd1 vccd1 _27377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_760 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24589_ _24589_/A vssd1 vssd1 vccd1 vccd1 _24598_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_156_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17130_ _17252_/A vssd1 vssd1 vccd1 vccd1 _17130_/X sky130_fd_sc_hd__clkbuf_2
X_14342_ _14342_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _14342_/Y sky130_fd_sc_hd__nor2_1
X_26328_ _20461_/X _26328_/D vssd1 vssd1 vccd1 vccd1 _26328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17061_ _17061_/A vssd1 vssd1 vccd1 vccd1 _17385_/S sky130_fd_sc_hd__buf_2
X_14273_ _26703_/Q _14270_/X _14271_/X _14272_/Y vssd1 vssd1 vccd1 vccd1 _26703_/D
+ sky130_fd_sc_hd__a31o_1
X_26259_ _20215_/X _26259_/D vssd1 vssd1 vccd1 vccd1 _26259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16012_ _27265_/Q _16012_/B vssd1 vssd1 vccd1 vccd1 _16030_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13224_ _13224_/A vssd1 vssd1 vccd1 vccd1 _27037_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _16249_/A vssd1 vssd1 vccd1 vccd1 _14766_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17963_ _17830_/X _17962_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _17963_/X sky130_fd_sc_hd__o21a_1
X_13086_ _14727_/A vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__buf_2
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19702_ _19694_/X _19695_/X _19696_/X _19697_/X _19698_/X _19699_/X vssd1 vssd1 vccd1
+ vccd1 _19703_/A sky130_fd_sc_hd__mux4_1
X_16914_ _16638_/A _16638_/B _16584_/Y vssd1 vssd1 vccd1 vccd1 _16915_/B sky130_fd_sc_hd__a21oi_1
XFILLER_26_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater407 _26047_/CLK vssd1 vssd1 vccd1 vccd1 _27356_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater418 _27327_/CLK vssd1 vssd1 vccd1 vccd1 _25958_/CLK sky130_fd_sc_hd__clkbuf_1
X_17894_ _18384_/A vssd1 vssd1 vccd1 vccd1 _17894_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater429 _26059_/CLK vssd1 vssd1 vccd1 vccd1 _26053_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19633_ _19621_/X _19622_/X _19623_/X _19624_/X _19625_/X _19626_/X vssd1 vssd1 vccd1
+ vccd1 _19634_/A sky130_fd_sc_hd__mux4_1
X_16845_ _16845_/A _16845_/B vssd1 vssd1 vccd1 vccd1 _16845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16776_ _16776_/A _16776_/B vssd1 vssd1 vccd1 vccd1 _16844_/B sky130_fd_sc_hd__or2_1
X_19564_ _26553_/Q _26521_/Q _26489_/Q _27065_/Q _18896_/X _18898_/X vssd1 vssd1 vccd1
+ vccd1 _19564_/X sky130_fd_sc_hd__mux4_1
X_13988_ _16536_/A vssd1 vssd1 vccd1 vccd1 _14361_/A sky130_fd_sc_hd__buf_2
XFILLER_20_1156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18515_ _26710_/Q _26678_/Q _26646_/Q _26614_/Q _17782_/X _17785_/X vssd1 vssd1 vccd1
+ vccd1 _18516_/A sky130_fd_sc_hd__mux4_2
X_15727_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15727_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _25075_/A vssd1 vssd1 vccd1 vccd1 _25297_/A sky130_fd_sc_hd__buf_4
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _19567_/A _19495_/B _19495_/C vssd1 vssd1 vccd1 vccd1 _19496_/A sky130_fd_sc_hd__and3_1
XFILLER_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15658_ _15680_/A vssd1 vssd1 vccd1 vccd1 _15667_/S sky130_fd_sc_hd__clkbuf_2
X_18446_ _18446_/A vssd1 vssd1 vccd1 vccd1 _25968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14609_ _26591_/Q _14602_/X _14605_/X _14608_/Y vssd1 vssd1 vccd1 vccd1 _26591_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18377_ _26960_/Q _26928_/Q _26896_/Q _26864_/Q _18244_/X _18269_/X vssd1 vssd1 vccd1
+ vccd1 _18377_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _26185_/Q _16252_/A _15595_/S vssd1 vssd1 vccd1 vccd1 _15590_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17328_ _25938_/Q _26004_/Q _17370_/S vssd1 vssd1 vccd1 vccd1 _17329_/B sky130_fd_sc_hd__mux2_1
XFILLER_193_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17259_ _27086_/Q _27118_/Q _17295_/S vssd1 vssd1 vccd1 vccd1 _17259_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20270_ _20270_/A vssd1 vssd1 vccd1 vccd1 _20336_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23960_ _27847_/Q _27151_/Q _25896_/Q _25864_/Q _23920_/X _23944_/X vssd1 vssd1 vccd1
+ vccd1 _23960_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22911_ _22943_/A vssd1 vssd1 vccd1 vccd1 _22911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23891_ _23889_/X _23890_/X _23891_/S vssd1 vssd1 vccd1 vccd1 _23891_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25630_ _25630_/A vssd1 vssd1 vccd1 vccd1 _25630_/X sky130_fd_sc_hd__clkbuf_1
X_22842_ _22858_/A vssd1 vssd1 vccd1 vccd1 _22842_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_519 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25561_ _25547_/X _25552_/X _25553_/X _24923_/B _25554_/X vssd1 vssd1 vccd1 vccd1
+ _25561_/X sky130_fd_sc_hd__o311a_1
X_22773_ _22767_/X _22768_/X _22769_/X _22770_/X _22771_/X _22772_/X vssd1 vssd1 vccd1
+ vccd1 _22774_/A sky130_fd_sc_hd__mux4_1
XFILLER_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27300_ _27686_/CLK _27300_/D vssd1 vssd1 vccd1 vccd1 _27300_/Q sky130_fd_sc_hd__dfxtp_1
X_24512_ _24589_/A vssd1 vssd1 vccd1 vccd1 _24554_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21724_ _21740_/A vssd1 vssd1 vccd1 vccd1 _21724_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25492_ _25552_/A vssd1 vssd1 vccd1 vccd1 _25492_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27231_ _27232_/CLK _27231_/D vssd1 vssd1 vccd1 vccd1 _27231_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24443_ _27620_/Q _24445_/B vssd1 vssd1 vccd1 vccd1 _24444_/A sky130_fd_sc_hd__and2_1
X_21655_ _21647_/X _21648_/X _21649_/X _21650_/X _21652_/X _21654_/X vssd1 vssd1 vccd1
+ vccd1 _21656_/A sky130_fd_sc_hd__mux4_1
XFILLER_200_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20606_ _20598_/X _20599_/X _20600_/X _20601_/X _20603_/X _20605_/X vssd1 vssd1 vccd1
+ vccd1 _20607_/A sky130_fd_sc_hd__mux4_1
X_27162_ _27541_/CLK _27162_/D vssd1 vssd1 vccd1 vccd1 _27162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24374_ _27569_/Q _24380_/B vssd1 vssd1 vccd1 vccd1 _24375_/A sky130_fd_sc_hd__and2_1
X_21586_ _21650_/A vssd1 vssd1 vccd1 vccd1 _21586_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26113_ _19707_/X _26113_/D vssd1 vssd1 vccd1 vccd1 _26113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23325_ _23325_/A _23325_/B _23325_/C vssd1 vssd1 vccd1 vccd1 _23332_/B sky130_fd_sc_hd__or3_1
XFILLER_192_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27093_ _27125_/CLK _27093_/D vssd1 vssd1 vccd1 vccd1 _27093_/Q sky130_fd_sc_hd__dfxtp_1
X_20537_ _20601_/A vssd1 vssd1 vccd1 vccd1 _20537_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_604 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26044_ _27358_/CLK _26044_/D vssd1 vssd1 vccd1 vccd1 _26044_/Q sky130_fd_sc_hd__dfxtp_1
X_20468_ _20500_/A vssd1 vssd1 vccd1 vccd1 _20468_/X sky130_fd_sc_hd__clkbuf_2
X_23256_ _27739_/Q vssd1 vssd1 vccd1 vccd1 _23256_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22207_ _22194_/X _22196_/X _22198_/X _22200_/X _22201_/X _22202_/X vssd1 vssd1 vccd1
+ vccd1 _22208_/A sky130_fd_sc_hd__mux4_1
XFILLER_161_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20399_ _20399_/A vssd1 vssd1 vccd1 vccd1 _20399_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23187_ _17428_/X _27131_/Q _23193_/S vssd1 vssd1 vccd1 vccd1 _23188_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22138_ _22138_/A vssd1 vssd1 vccd1 vccd1 _22138_/X sky130_fd_sc_hd__clkbuf_1
X_27995_ _27995_/A _15886_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_854 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26946_ _22622_/X _26946_/D vssd1 vssd1 vccd1 vccd1 _26946_/Q sky130_fd_sc_hd__dfxtp_1
X_14960_ _15043_/B vssd1 vssd1 vccd1 vccd1 _14960_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22069_ _22085_/A vssd1 vssd1 vccd1 vccd1 _22069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13911_ _26822_/Q _13906_/X _13899_/X _13910_/Y vssd1 vssd1 vccd1 vccd1 _26822_/D
+ sky130_fd_sc_hd__a31o_1
X_26877_ _22380_/X _26877_/D vssd1 vssd1 vccd1 vccd1 _26877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14891_ _14891_/A vssd1 vssd1 vccd1 vccd1 _26488_/D sky130_fd_sc_hd__clkbuf_1
X_16630_ _16664_/A _16664_/B _16629_/X vssd1 vssd1 vccd1 vccd1 _16631_/B sky130_fd_sc_hd__a21oi_1
X_13842_ _13936_/A _13847_/B vssd1 vssd1 vccd1 vccd1 _13842_/Y sky130_fd_sc_hd__nor2_1
X_25828_ _25996_/CLK _25828_/D vssd1 vssd1 vccd1 vccd1 _25828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16561_ _16561_/A _16561_/B vssd1 vssd1 vccd1 vccd1 _16570_/B sky130_fd_sc_hd__xor2_1
X_13773_ _13827_/A vssd1 vssd1 vccd1 vccd1 _13785_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25759_ _25805_/S vssd1 vssd1 vccd1 vccd1 _25768_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15512_ _13139_/X _26219_/Q _15512_/S vssd1 vssd1 vccd1 vccd1 _15513_/A sky130_fd_sc_hd__mux2_1
X_18300_ _18300_/A _18207_/X vssd1 vssd1 vccd1 vccd1 _18300_/X sky130_fd_sc_hd__or2b_1
X_19280_ _19438_/A vssd1 vssd1 vccd1 vccd1 _19419_/A sky130_fd_sc_hd__clkbuf_1
X_16492_ _16493_/B _16493_/C _16809_/B vssd1 vssd1 vccd1 vccd1 _16494_/A sky130_fd_sc_hd__a21oi_1
XFILLER_71_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18231_ _26281_/Q _26249_/Q _26217_/Q _26185_/Q _18185_/X _18209_/X vssd1 vssd1 vccd1
+ vccd1 _18231_/X sky130_fd_sc_hd__mux4_1
XFILLER_176_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27429_ _27437_/CLK _27429_/D vssd1 vssd1 vccd1 vccd1 _27429_/Q sky130_fd_sc_hd__dfxtp_1
X_15443_ _26250_/Q _13369_/X _15451_/S vssd1 vssd1 vccd1 vccd1 _15444_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18162_ _18437_/A vssd1 vssd1 vccd1 vccd1 _18162_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15374_ _15374_/A vssd1 vssd1 vccd1 vccd1 _26281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17113_ _17111_/X _17112_/X _17113_/S vssd1 vssd1 vccd1 vccd1 _17113_/X sky130_fd_sc_hd__mux2_1
X_14325_ _14412_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18093_ _18093_/A _17799_/X vssd1 vssd1 vccd1 vccd1 _18093_/X sky130_fd_sc_hd__or2b_1
XFILLER_8_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ _25814_/Q _26013_/Q _17097_/S vssd1 vssd1 vccd1 vccd1 _17044_/X sky130_fd_sc_hd__mux2_1
X_14256_ _14296_/A vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13207_ _13207_/A vssd1 vssd1 vccd1 vccd1 _27040_/D sky130_fd_sc_hd__clkbuf_1
X_14187_ _14363_/A _14187_/B vssd1 vssd1 vccd1 vccd1 _14187_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_800 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _16271_/A vssd1 vssd1 vccd1 vccd1 _14756_/A sky130_fd_sc_hd__clkbuf_4
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _19113_/A _18995_/B vssd1 vssd1 vccd1 vccd1 _18995_/X sky130_fd_sc_hd__or2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _17936_/X _17941_/X _17945_/X _17854_/X _17856_/X vssd1 vssd1 vccd1 vccd1
+ _17947_/C sky130_fd_sc_hd__a221o_1
X_13069_ _13069_/A vssd1 vssd1 vccd1 vccd1 _27063_/D sky130_fd_sc_hd__clkbuf_1
Xrepeater204 _25884_/CLK vssd1 vssd1 vccd1 vccd1 _27835_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater215 _27790_/CLK vssd1 vssd1 vccd1 vccd1 _27232_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater226 _25974_/CLK vssd1 vssd1 vccd1 vccd1 _26065_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater237 _27751_/CLK vssd1 vssd1 vccd1 vccd1 _27729_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater248 _27527_/CLK vssd1 vssd1 vccd1 vccd1 _27726_/CLK sky130_fd_sc_hd__clkbuf_1
X_17877_ _18305_/A vssd1 vssd1 vccd1 vccd1 _17877_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater259 _27611_/CLK vssd1 vssd1 vccd1 vccd1 _27612_/CLK sky130_fd_sc_hd__clkbuf_1
X_19616_ _19616_/A vssd1 vssd1 vccd1 vccd1 _19616_/X sky130_fd_sc_hd__clkbuf_1
X_16828_ _16821_/Y _16827_/Y _16812_/A vssd1 vssd1 vccd1 vccd1 _16841_/B sky130_fd_sc_hd__o21a_1
XFILLER_93_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19547_ _19545_/X _19546_/X _19565_/S vssd1 vssd1 vccd1 vccd1 _19547_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16759_ _16759_/A _16759_/B vssd1 vssd1 vccd1 vccd1 _16842_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19478_ _26965_/Q _26933_/Q _26901_/Q _26869_/Q _18824_/X _19412_/X vssd1 vssd1 vccd1
+ vccd1 _19478_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18429_ _18426_/X _18428_/X _18532_/S vssd1 vssd1 vccd1 vccd1 _18429_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21440_ _21440_/A vssd1 vssd1 vccd1 vccd1 _21440_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21371_ _21357_/X _21358_/X _21359_/X _21360_/X _21361_/X _21362_/X vssd1 vssd1 vccd1
+ vccd1 _21372_/A sky130_fd_sc_hd__mux4_1
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23110_ _27375_/Q _24002_/A vssd1 vssd1 vccd1 vccd1 _23167_/A sky130_fd_sc_hd__and2_1
X_20322_ _20322_/A vssd1 vssd1 vccd1 vccd1 _20322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24090_ _24090_/A vssd1 vssd1 vccd1 vccd1 _27320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_446 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20253_ _20322_/A vssd1 vssd1 vccd1 vccd1 _20253_/X sky130_fd_sc_hd__clkbuf_2
X_23041_ _23041_/A vssd1 vssd1 vccd1 vccd1 _27066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20184_ _20270_/A vssd1 vssd1 vccd1 vccd1 _20250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26800_ _22116_/X _26800_/D vssd1 vssd1 vccd1 vccd1 _26800_/Q sky130_fd_sc_hd__dfxtp_1
X_27780_ _27781_/CLK _27780_/D vssd1 vssd1 vccd1 vccd1 _27780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24992_ _27828_/Q _27132_/Q _25877_/Q _25845_/Q _24972_/X _24991_/X vssd1 vssd1 vccd1
+ vccd1 _24992_/X sky130_fd_sc_hd__mux4_1
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26731_ _21872_/X _26731_/D vssd1 vssd1 vccd1 vccd1 _26731_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23943_ _23990_/A vssd1 vssd1 vccd1 vccd1 _23943_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26662_ _21626_/X _26662_/D vssd1 vssd1 vccd1 vccd1 _26662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23874_ _27838_/Q _27142_/Q _25887_/Q _25855_/Q _23873_/X _23850_/X vssd1 vssd1 vccd1
+ vccd1 _23874_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25613_ _25560_/X _25356_/B _25612_/X _25543_/X vssd1 vssd1 vccd1 vccd1 _25613_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22825_ _22857_/A vssd1 vssd1 vccd1 vccd1 _22825_/X sky130_fd_sc_hd__clkbuf_2
X_26593_ _21386_/X _26593_/D vssd1 vssd1 vccd1 vccd1 _26593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25544_ _25530_/X _25253_/B _25542_/X _25543_/X vssd1 vssd1 vccd1 vccd1 _25544_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22756_ _22772_/A vssd1 vssd1 vccd1 vccd1 _22756_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21707_ _21739_/A vssd1 vssd1 vccd1 vccd1 _21707_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25475_ _27696_/Q _25448_/X _25449_/X vssd1 vssd1 vccd1 vccd1 _25475_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22687_ _22681_/X _22682_/X _22683_/X _22684_/X _22685_/X _22686_/X vssd1 vssd1 vccd1
+ vccd1 _22688_/A sky130_fd_sc_hd__mux4_1
XFILLER_13_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27214_ _27214_/CLK _27214_/D vssd1 vssd1 vccd1 vccd1 _27214_/Q sky130_fd_sc_hd__dfxtp_1
X_24426_ _24426_/A vssd1 vssd1 vccd1 vccd1 _27491_/D sky130_fd_sc_hd__clkbuf_1
X_21638_ _21638_/A vssd1 vssd1 vccd1 vccd1 _21638_/X sky130_fd_sc_hd__clkbuf_1
X_27145_ _27145_/CLK _27145_/D vssd1 vssd1 vccd1 vccd1 _27145_/Q sky130_fd_sc_hd__dfxtp_1
X_24357_ _27561_/Q _24361_/B vssd1 vssd1 vccd1 vccd1 _24358_/A sky130_fd_sc_hd__and2_1
X_21569_ _21561_/X _21562_/X _21563_/X _21564_/X _21566_/X _21568_/X vssd1 vssd1 vccd1
+ vccd1 _21570_/A sky130_fd_sc_hd__mux4_1
XFILLER_181_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14110_ _14374_/A _14112_/B vssd1 vssd1 vccd1 vccd1 _14110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23308_ _27730_/Q _23305_/Y _23302_/Y input64/X _23307_/X vssd1 vssd1 vccd1 vccd1
+ _23309_/C sky130_fd_sc_hd__a221o_1
X_27076_ _27076_/CLK _27076_/D vssd1 vssd1 vccd1 vccd1 _27076_/Q sky130_fd_sc_hd__dfxtp_1
X_15090_ _14772_/X _26406_/Q _15090_/S vssd1 vssd1 vccd1 vccd1 _15091_/A sky130_fd_sc_hd__mux2_1
X_24288_ _24288_/A vssd1 vssd1 vccd1 vccd1 _27422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ _26784_/Q _14024_/X _14038_/X _14040_/Y vssd1 vssd1 vccd1 vccd1 _26784_/D
+ sky130_fd_sc_hd__a31o_1
X_26027_ _27083_/CLK _26027_/D vssd1 vssd1 vccd1 vccd1 _26027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23239_ _23239_/A vssd1 vssd1 vccd1 vccd1 _23248_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_181_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27954__440 vssd1 vssd1 vccd1 vccd1 _27954__440/HI _27954_/A sky130_fd_sc_hd__conb_1
XFILLER_4_489 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17800_ _18360_/A vssd1 vssd1 vccd1 vccd1 _18085_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15992_ _15992_/A vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__clkbuf_1
X_18780_ _18897_/A vssd1 vssd1 vccd1 vccd1 _18923_/A sky130_fd_sc_hd__clkbuf_2
X_27978_ _27978_/A _15906_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
XFILLER_122_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_600 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17731_ _27425_/Q vssd1 vssd1 vccd1 vccd1 _17731_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14943_ _14791_/X _26464_/Q _14951_/S vssd1 vssd1 vccd1 vccd1 _14944_/A sky130_fd_sc_hd__mux2_1
X_26929_ _22560_/X _26929_/D vssd1 vssd1 vccd1 vccd1 _26929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_603 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17662_ _17662_/A vssd1 vssd1 vccd1 vccd1 _25901_/D sky130_fd_sc_hd__clkbuf_1
X_14874_ _14874_/A vssd1 vssd1 vccd1 vccd1 _26495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ _19401_/A vssd1 vssd1 vccd1 vccd1 _19401_/X sky130_fd_sc_hd__buf_2
XFILLER_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13825_ _13917_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13825_/Y sky130_fd_sc_hd__nor2_1
X_16613_ _16093_/X _16610_/X _16611_/X _16612_/X vssd1 vssd1 vccd1 vccd1 _24240_/A
+ sky130_fd_sc_hd__a22o_1
X_17593_ _17514_/X _25871_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17594_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16544_ _16815_/B _16545_/B _16666_/B _16629_/B vssd1 vssd1 vccd1 vccd1 _16544_/X
+ sky130_fd_sc_hd__o211a_1
X_19332_ _26414_/Q _26382_/Q _26350_/Q _26318_/Q _19331_/X _19240_/X vssd1 vssd1 vccd1
+ vccd1 _19332_/X sky130_fd_sc_hd__mux4_1
X_13756_ _26876_/Q _13750_/X _13745_/X _13755_/Y vssd1 vssd1 vccd1 vccd1 _26876_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19263_ _19191_/X _19262_/X _19194_/X vssd1 vssd1 vccd1 vccd1 _19263_/X sky130_fd_sc_hd__o21a_1
X_16475_ _16479_/A _16479_/B vssd1 vssd1 vccd1 vccd1 _16475_/Y sky130_fd_sc_hd__nor2_1
X_13687_ _13868_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13687_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18214_ _18486_/A vssd1 vssd1 vccd1 vccd1 _18214_/X sky130_fd_sc_hd__clkbuf_2
X_15426_ _15426_/A vssd1 vssd1 vccd1 vccd1 _26258_/D sky130_fd_sc_hd__clkbuf_1
X_19194_ _19488_/A vssd1 vssd1 vccd1 vccd1 _19194_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15357_ _14740_/X _26288_/Q _15357_/S vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__mux2_1
X_18145_ _18138_/X _18140_/X _18144_/X _18026_/X _18122_/X vssd1 vssd1 vccd1 vccd1
+ _18146_/C sky130_fd_sc_hd__a221o_1
XFILLER_102_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_881 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ _26689_/Q _14296_/X _14297_/X _14307_/Y vssd1 vssd1 vccd1 vccd1 _26689_/D
+ sky130_fd_sc_hd__a31o_1
X_18076_ _18067_/X _18071_/X _18075_/X _18026_/X _17990_/X vssd1 vssd1 vccd1 vccd1
+ _18077_/C sky130_fd_sc_hd__a221o_1
X_15288_ _15288_/A vssd1 vssd1 vccd1 vccd1 _26319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17027_ _17027_/A vssd1 vssd1 vccd1 vccd1 _27917_/A sky130_fd_sc_hd__clkbuf_1
X_14239_ _15695_/A _15695_/B _15695_/C vssd1 vssd1 vccd1 vccd1 _14534_/B sky130_fd_sc_hd__and3b_2
XFILLER_171_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_660 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18978_ _26143_/Q _26079_/Q _27007_/Q _26975_/Q _18882_/X _18950_/X vssd1 vssd1 vccd1
+ vccd1 _18979_/B sky130_fd_sc_hd__mux4_1
XFILLER_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17929_ _26685_/Q _26653_/Q _26621_/Q _26589_/Q _17865_/X _17928_/X vssd1 vssd1 vccd1
+ vccd1 _17930_/A sky130_fd_sc_hd__mux4_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20940_ _20956_/A vssd1 vssd1 vccd1 vccd1 _20940_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20871_ input3/X vssd1 vssd1 vccd1 vccd1 _22616_/A sky130_fd_sc_hd__buf_6
XFILLER_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22610_ _22610_/A vssd1 vssd1 vccd1 vccd1 _22610_/X sky130_fd_sc_hd__clkbuf_1
X_23590_ _23590_/A vssd1 vssd1 vccd1 vccd1 _27217_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22541_ _22889_/A vssd1 vssd1 vccd1 vccd1 _22610_/A sky130_fd_sc_hd__buf_2
XFILLER_22_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25260_ _25265_/B _25260_/B vssd1 vssd1 vccd1 vccd1 _25261_/B sky130_fd_sc_hd__xor2_1
XFILLER_72_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22472_ _22520_/A vssd1 vssd1 vccd1 vccd1 _22472_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24211_ _24363_/A vssd1 vssd1 vccd1 vccd1 _24380_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_194_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21423_ _21408_/X _21410_/X _21412_/X _21414_/X _21415_/X _21416_/X vssd1 vssd1 vccd1
+ vccd1 _21424_/A sky130_fd_sc_hd__mux4_1
XFILLER_182_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25191_ _25191_/A _25191_/B vssd1 vssd1 vccd1 vccd1 _25192_/B sky130_fd_sc_hd__xnor2_1
XFILLER_33_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24142_ _24175_/A vssd1 vssd1 vccd1 vccd1 _24151_/B sky130_fd_sc_hd__clkbuf_1
X_21354_ _21354_/A vssd1 vssd1 vccd1 vccd1 _21354_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20305_ _20337_/A vssd1 vssd1 vccd1 vccd1 _20305_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24073_ _24073_/A vssd1 vssd1 vccd1 vccd1 _27313_/D sky130_fd_sc_hd__clkbuf_1
X_21285_ _21301_/A vssd1 vssd1 vccd1 vccd1 _21285_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_522 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23024_ _23024_/A vssd1 vssd1 vccd1 vccd1 _23024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20236_ _20236_/A vssd1 vssd1 vccd1 vccd1 _20236_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20167_ _20236_/A vssd1 vssd1 vccd1 vccd1 _20167_/X sky130_fd_sc_hd__clkbuf_2
X_27832_ _27832_/CLK _27832_/D vssd1 vssd1 vccd1 vccd1 _27832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24975_ _25035_/A vssd1 vssd1 vccd1 vccd1 _24975_/X sky130_fd_sc_hd__buf_2
X_27763_ _27766_/CLK _27763_/D vssd1 vssd1 vccd1 vccd1 _27763_/Q sky130_fd_sc_hd__dfxtp_2
X_20098_ _20270_/A vssd1 vssd1 vccd1 vccd1 _20164_/A sky130_fd_sc_hd__buf_2
XFILLER_188_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23926_ _27083_/Q _23907_/X _23908_/X _27115_/Q _23909_/X vssd1 vssd1 vccd1 vccd1
+ _23926_/X sky130_fd_sc_hd__a221o_1
X_26714_ _21808_/X _26714_/D vssd1 vssd1 vccd1 vccd1 _26714_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27694_ _27695_/CLK _27694_/D vssd1 vssd1 vccd1 vccd1 _27694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_636 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26645_ _21570_/X _26645_/D vssd1 vssd1 vccd1 vccd1 _26645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23857_ _27076_/Q _27108_/Q _23892_/S vssd1 vssd1 vccd1 vccd1 _23857_/X sky130_fd_sc_hd__mux2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _13649_/A vssd1 vssd1 vccd1 vccd1 _13621_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22808_ _22872_/A vssd1 vssd1 vccd1 vccd1 _22808_/X sky130_fd_sc_hd__clkbuf_1
X_14590_ _15751_/A _14597_/B vssd1 vssd1 vccd1 vccd1 _14590_/Y sky130_fd_sc_hd__nor2_1
X_26576_ _21334_/X _26576_/D vssd1 vssd1 vccd1 vccd1 _26576_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23788_ _23785_/X _23787_/X _23795_/S vssd1 vssd1 vccd1 vccd1 _23788_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13541_ _14500_/A vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__clkbuf_2
X_25527_ _25592_/A vssd1 vssd1 vccd1 vccd1 _25527_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22739_ _22771_/A vssd1 vssd1 vccd1 vccd1 _22739_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16260_ _26061_/Q _16137_/X _16138_/Y _13127_/A vssd1 vssd1 vccd1 vccd1 _16260_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _26962_/Q _13464_/X _13457_/X _13471_/Y vssd1 vssd1 vccd1 vccd1 _26962_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25458_ _25438_/X _25139_/B _25457_/X _25452_/X vssd1 vssd1 vccd1 vccd1 _25458_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _15211_/A vssd1 vssd1 vccd1 vccd1 _26353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24409_ _27585_/Q _24411_/B vssd1 vssd1 vccd1 vccd1 _24410_/A sky130_fd_sc_hd__and2_1
X_16191_ _16191_/A _16191_/B _16197_/C vssd1 vssd1 vccd1 vccd1 _16191_/X sky130_fd_sc_hd__and3_1
X_25389_ _27734_/Q input45/X _25391_/S vssd1 vssd1 vccd1 vccd1 _25390_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27128_ _27674_/CLK _27128_/D vssd1 vssd1 vccd1 vccd1 _27128_/Q sky130_fd_sc_hd__dfxtp_1
X_15142_ _15188_/S vssd1 vssd1 vccd1 vccd1 _15151_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_153_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19950_ _19940_/X _19941_/X _19942_/X _19943_/X _19944_/X _19945_/X vssd1 vssd1 vccd1
+ vccd1 _19951_/A sky130_fd_sc_hd__mux4_1
X_15073_ _14747_/X _26414_/Q _15079_/S vssd1 vssd1 vccd1 vccd1 _15074_/A sky130_fd_sc_hd__mux2_1
X_27059_ _23008_/X _27059_/D vssd1 vssd1 vccd1 vccd1 _27059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _14090_/A vssd1 vssd1 vccd1 vccd1 _14024_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18901_ _18923_/A vssd1 vssd1 vccd1 vccd1 _18901_/X sky130_fd_sc_hd__buf_4
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19881_ _19881_/A vssd1 vssd1 vccd1 vccd1 _19881_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18832_ _26522_/Q _26490_/Q _26458_/Q _27034_/Q _18829_/X _18831_/X vssd1 vssd1 vccd1
+ vccd1 _18832_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18763_ _27600_/Q vssd1 vssd1 vccd1 vccd1 _19428_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15975_ _15979_/A vssd1 vssd1 vccd1 vccd1 _15975_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17714_ _17714_/A vssd1 vssd1 vccd1 vccd1 _25923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14926_ _14926_/A vssd1 vssd1 vccd1 vccd1 _26472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18694_ _26010_/Q _17673_/X _18702_/S vssd1 vssd1 vccd1 vccd1 _18695_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17645_ _17485_/X _25894_/Q _17645_/S vssd1 vssd1 vccd1 vccd1 _17646_/A sky130_fd_sc_hd__mux2_1
X_14857_ _26502_/Q _13382_/X _14857_/S vssd1 vssd1 vccd1 vccd1 _14858_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ _13900_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13808_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17576_ _17488_/X _25863_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17577_/A sky130_fd_sc_hd__mux2_1
X_14788_ _16206_/A vssd1 vssd1 vccd1 vccd1 _14788_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19315_ _26830_/Q _26798_/Q _26766_/Q _26734_/Q _19203_/X _19248_/X vssd1 vssd1 vccd1
+ vccd1 _19316_/B sky130_fd_sc_hd__mux4_1
XFILLER_182_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13739_ _26883_/Q _13737_/X _13732_/X _13738_/Y vssd1 vssd1 vccd1 vccd1 _26883_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16527_ _16908_/A _16552_/B vssd1 vssd1 vccd1 vccd1 _16911_/A sky130_fd_sc_hd__xnor2_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19246_ _19362_/A _19246_/B _19246_/C vssd1 vssd1 vccd1 vccd1 _19247_/A sky130_fd_sc_hd__and3_1
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16458_ _14766_/A _16384_/A _16374_/A _25958_/Q _16457_/X vssd1 vssd1 vccd1 vccd1
+ _16470_/A sky130_fd_sc_hd__a221o_2
XFILLER_104_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15409_ _15477_/S vssd1 vssd1 vccd1 vccd1 _15418_/S sky130_fd_sc_hd__clkbuf_2
X_19177_ _26824_/Q _26792_/Q _26760_/Q _26728_/Q _19039_/X _19111_/X vssd1 vssd1 vccd1
+ vccd1 _19178_/B sky130_fd_sc_hd__mux4_1
XFILLER_176_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16389_ _16447_/B _16357_/A _16745_/A _16369_/X vssd1 vssd1 vccd1 vccd1 _16390_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18128_ _18455_/A vssd1 vssd1 vccd1 vccd1 _18427_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_184_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18059_ _26818_/Q _26786_/Q _26754_/Q _26722_/Q _18034_/X _18058_/X vssd1 vssd1 vccd1
+ vccd1 _18059_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21070_ _21070_/A vssd1 vssd1 vccd1 vccd1 _21070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20021_ _20021_/A vssd1 vssd1 vccd1 vccd1 _20021_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24760_ _24801_/A vssd1 vssd1 vccd1 vccd1 _24760_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21972_ _21972_/A vssd1 vssd1 vccd1 vccd1 _21972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23711_ _23711_/A vssd1 vssd1 vccd1 vccd1 _27259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20923_ _20955_/A vssd1 vssd1 vccd1 vccd1 _20923_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24691_ _24386_/A _24687_/X _24689_/X _24690_/X vssd1 vssd1 vccd1 vccd1 _27593_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26430_ _20823_/X _26430_/D vssd1 vssd1 vccd1 vccd1 _26430_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23642_ _27231_/Q vssd1 vssd1 vccd1 vccd1 _25003_/S sky130_fd_sc_hd__clkbuf_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20854_ _20848_/X _20849_/X _20850_/X _20851_/X _20852_/X _20853_/X vssd1 vssd1 vccd1
+ vccd1 _20855_/A sky130_fd_sc_hd__mux4_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26361_ _20575_/X _26361_/D vssd1 vssd1 vccd1 vccd1 _26361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23573_ _24906_/A _27213_/Q _23576_/S vssd1 vssd1 vccd1 vccd1 _23574_/B sky130_fd_sc_hd__mux2_1
X_20785_ _20785_/A vssd1 vssd1 vccd1 vccd1 _20785_/X sky130_fd_sc_hd__clkbuf_1
X_25312_ _25329_/C _25312_/B vssd1 vssd1 vccd1 vccd1 _25313_/B sky130_fd_sc_hd__xnor2_1
X_22524_ _22597_/A vssd1 vssd1 vccd1 vccd1 _22524_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26292_ _20329_/X _26292_/D vssd1 vssd1 vccd1 vccd1 _26292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25243_ _25250_/A _25243_/B vssd1 vssd1 vccd1 vccd1 _25244_/B sky130_fd_sc_hd__nor2_1
X_22455_ _22455_/A vssd1 vssd1 vccd1 vccd1 _22521_/A sky130_fd_sc_hd__buf_2
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21406_ _21406_/A vssd1 vssd1 vccd1 vccd1 _21406_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25174_ _25182_/A _25174_/B vssd1 vssd1 vccd1 vccd1 _25174_/Y sky130_fd_sc_hd__nand2_1
X_22386_ _22434_/A vssd1 vssd1 vccd1 vccd1 _22386_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_850 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24125_ _24125_/A vssd1 vssd1 vccd1 vccd1 _27336_/D sky130_fd_sc_hd__clkbuf_1
X_21337_ _21322_/X _21324_/X _21326_/X _21328_/X _21329_/X _21330_/X vssd1 vssd1 vccd1
+ vccd1 _21338_/A sky130_fd_sc_hd__mux4_1
XFILLER_135_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1078 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24056_ _24056_/A vssd1 vssd1 vccd1 vccd1 _27305_/D sky130_fd_sc_hd__clkbuf_1
X_21268_ _21268_/A vssd1 vssd1 vccd1 vccd1 _21268_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23007_ _22993_/X _22994_/X _22995_/X _22996_/X _22997_/X _22998_/X vssd1 vssd1 vccd1
+ vccd1 _23008_/A sky130_fd_sc_hd__mux4_1
XFILLER_104_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20219_ _20251_/A vssd1 vssd1 vccd1 vccd1 _20219_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21199_ _21199_/A vssd1 vssd1 vccd1 vccd1 _21199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27815_ _25702_/X _27815_/D vssd1 vssd1 vccd1 vccd1 _27815_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _24980_/S vssd1 vssd1 vccd1 vccd1 _15760_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _27811_/Q _12976_/B vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__and2_1
X_27746_ _27746_/CLK _27746_/D vssd1 vssd1 vccd1 vccd1 _27746_/Q sky130_fd_sc_hd__dfxtp_1
X_24958_ _27668_/Q _24935_/X _24957_/Y _24938_/X vssd1 vssd1 vccd1 vccd1 _27668_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14792_/A vssd1 vssd1 vccd1 vccd1 _14811_/S sky130_fd_sc_hd__buf_2
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23909_ _24003_/A vssd1 vssd1 vccd1 vccd1 _23909_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15691_ _13234_/X _26139_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15692_/A sky130_fd_sc_hd__mux2_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24889_ _24889_/A _24889_/B vssd1 vssd1 vccd1 vccd1 _24889_/Y sky130_fd_sc_hd__nand2_1
X_27677_ _27677_/CLK _27677_/D vssd1 vssd1 vccd1 vccd1 _27968_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _26580_/Q _14630_/X _14640_/X _14641_/Y vssd1 vssd1 vccd1 vccd1 _26580_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17430_ _17430_/A vssd1 vssd1 vccd1 vccd1 _25812_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26628_ _21510_/X _26628_/D vssd1 vssd1 vccd1 vccd1 _26628_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14573_ _14599_/A vssd1 vssd1 vccd1 vccd1 _14584_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17361_ _17338_/X _17361_/B vssd1 vssd1 vccd1 vccd1 _17361_/X sky130_fd_sc_hd__and2b_1
XFILLER_198_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26559_ _21268_/X _26559_/D vssd1 vssd1 vccd1 vccd1 _26559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19100_ _19399_/A vssd1 vssd1 vccd1 vccd1 _19100_/X sky130_fd_sc_hd__clkbuf_2
X_13524_ _27347_/Q _13021_/A _13102_/X _27315_/Q _13164_/X vssd1 vssd1 vccd1 vccd1
+ _16442_/A sky130_fd_sc_hd__a221oi_4
X_16312_ _16402_/A vssd1 vssd1 vccd1 vccd1 _16312_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17292_ _25834_/Q _26033_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19031_ _26401_/Q _26369_/Q _26337_/Q _26305_/Q _18887_/X _18982_/X vssd1 vssd1 vccd1
+ vccd1 _19031_/X sky130_fd_sc_hd__mux4_1
X_16243_ _16243_/A _16277_/B vssd1 vssd1 vccd1 vccd1 _16243_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ _26965_/Q _13435_/X _13429_/X _13454_/Y vssd1 vssd1 vccd1 vccd1 _26965_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_103_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16174_ _27377_/Q vssd1 vssd1 vccd1 vccd1 _16342_/A sky130_fd_sc_hd__inv_2
X_13386_ _13402_/A vssd1 vssd1 vccd1 vccd1 _13399_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_541 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15125_ _26391_/Q _13328_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15126_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19933_ _19933_/A vssd1 vssd1 vccd1 vccd1 _19933_/X sky130_fd_sc_hd__clkbuf_1
X_15056_ _15056_/A vssd1 vssd1 vccd1 vccd1 _26422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14007_ _14374_/A _14010_/B vssd1 vssd1 vccd1 vccd1 _14007_/Y sky130_fd_sc_hd__nor2_1
X_19864_ _19850_/X _19851_/X _19852_/X _19853_/X _19854_/X _19855_/X vssd1 vssd1 vccd1
+ vccd1 _19865_/A sky130_fd_sc_hd__mux4_1
XFILLER_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18815_ _18922_/A vssd1 vssd1 vccd1 vccd1 _19317_/A sky130_fd_sc_hd__clkbuf_4
X_19795_ _19795_/A vssd1 vssd1 vccd1 vccd1 _19795_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18746_ _26034_/Q _17753_/X _18746_/S vssd1 vssd1 vccd1 vccd1 _18747_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15958_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15958_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _14955_/S vssd1 vssd1 vccd1 vccd1 _14918_/S sky130_fd_sc_hd__clkbuf_2
X_18677_ _26003_/Q _17756_/X _18685_/S vssd1 vssd1 vccd1 vccd1 _18678_/A sky130_fd_sc_hd__mux2_1
X_15889_ _15893_/A vssd1 vssd1 vccd1 vccd1 _15889_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17628_ _17460_/X _25886_/Q _17634_/S vssd1 vssd1 vccd1 vccd1 _17629_/A sky130_fd_sc_hd__mux2_1
XFILLER_197_909 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ _17559_/A vssd1 vssd1 vccd1 vccd1 _25855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20570_ _20586_/A vssd1 vssd1 vccd1 vccd1 _20570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19229_ _19387_/A vssd1 vssd1 vccd1 vccd1 _19229_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22240_ _22240_/A vssd1 vssd1 vccd1 vccd1 _22240_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22171_ _22157_/X _22158_/X _22159_/X _22160_/X _22161_/X _22162_/X vssd1 vssd1 vccd1
+ vccd1 _22172_/A sky130_fd_sc_hd__mux4_1
XFILLER_172_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21122_ _21122_/A vssd1 vssd1 vccd1 vccd1 _21122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25930_ _25996_/CLK _25930_/D vssd1 vssd1 vccd1 vccd1 _25930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21053_ _21039_/X _21040_/X _21041_/X _21042_/X _21044_/X _21046_/X vssd1 vssd1 vccd1
+ vccd1 _21054_/A sky130_fd_sc_hd__mux4_1
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20004_ _19988_/X _19989_/X _19990_/X _19991_/X _19994_/X _19997_/X vssd1 vssd1 vccd1
+ vccd1 _20005_/A sky130_fd_sc_hd__mux4_1
XFILLER_101_633 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25861_ _27148_/CLK _25861_/D vssd1 vssd1 vccd1 vccd1 _25861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24812_ _27637_/Q _24798_/X _24811_/Y _24801_/X vssd1 vssd1 vccd1 vccd1 _27637_/D
+ sky130_fd_sc_hd__o211a_1
X_27600_ _27600_/CLK _27600_/D vssd1 vssd1 vccd1 vccd1 _27600_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25792_ _25792_/A vssd1 vssd1 vccd1 vccd1 _25801_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24743_ _24844_/A vssd1 vssd1 vccd1 vccd1 _24744_/A sky130_fd_sc_hd__inv_2
X_27531_ _27531_/CLK _27531_/D vssd1 vssd1 vccd1 vccd1 _27531_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21955_ _21949_/X _21950_/X _21951_/X _21952_/X _21953_/X _21954_/X vssd1 vssd1 vccd1
+ vccd1 _21956_/A sky130_fd_sc_hd__mux4_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27462_ _27462_/CLK _27462_/D vssd1 vssd1 vccd1 vccd1 _27462_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _20954_/A vssd1 vssd1 vccd1 vccd1 _20906_/X sky130_fd_sc_hd__clkbuf_1
X_24674_ _25540_/A vssd1 vssd1 vccd1 vccd1 _24685_/B sky130_fd_sc_hd__clkbuf_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21886_ _21886_/A vssd1 vssd1 vccd1 vccd1 _21886_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26413_ _20751_/X _26413_/D vssd1 vssd1 vccd1 vccd1 _26413_/Q sky130_fd_sc_hd__dfxtp_1
X_23625_ _23625_/A vssd1 vssd1 vccd1 vccd1 _27226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20837_ _20853_/A vssd1 vssd1 vccd1 vccd1 _20837_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27393_ _27394_/CLK _27393_/D vssd1 vssd1 vccd1 vccd1 _27393_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26344_ _20511_/X _26344_/D vssd1 vssd1 vccd1 vccd1 _26344_/Q sky130_fd_sc_hd__dfxtp_1
X_23556_ _27766_/Q _27208_/Q _23559_/S vssd1 vssd1 vccd1 vccd1 _23557_/B sky130_fd_sc_hd__mux2_1
XFILLER_196_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20768_ _20754_/X _20755_/X _20756_/X _20757_/X _20758_/X _20759_/X vssd1 vssd1 vccd1
+ vccd1 _20769_/A sky130_fd_sc_hd__mux4_1
XFILLER_196_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22507_ _22507_/A vssd1 vssd1 vccd1 vccd1 _22507_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26275_ _20277_/X _26275_/D vssd1 vssd1 vccd1 vccd1 _26275_/Q sky130_fd_sc_hd__dfxtp_1
X_23487_ _25132_/A vssd1 vssd1 vccd1 vccd1 _23487_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_20699_ _20699_/A vssd1 vssd1 vccd1 vccd1 _20699_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_28014_ _28014_/A _15977_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_25226_ _27534_/Q _27502_/Q vssd1 vssd1 vccd1 vccd1 _25228_/A sky130_fd_sc_hd__nand2_1
X_13240_ _14810_/A vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1129 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22438_ _22507_/A vssd1 vssd1 vccd1 vccd1 _22438_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25157_ _25157_/A _25157_/B vssd1 vssd1 vccd1 vccd1 _25158_/B sky130_fd_sc_hd__xnor2_1
X_13171_ _16157_/A vssd1 vssd1 vccd1 vccd1 _14775_/A sky130_fd_sc_hd__clkbuf_4
X_22369_ _22455_/A vssd1 vssd1 vccd1 vccd1 _22435_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24108_ _24119_/A vssd1 vssd1 vccd1 vccd1 _24117_/B sky130_fd_sc_hd__clkbuf_1
X_25088_ _27079_/Q _27111_/Q _25088_/S vssd1 vssd1 vccd1 vccd1 _25088_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24039_ _27096_/Q _27128_/Q _24046_/S vssd1 vssd1 vccd1 vccd1 _24039_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16930_ _27595_/Q _24208_/A _24209_/A _27596_/Q vssd1 vssd1 vccd1 vccd1 _16930_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16861_ _16738_/A _16858_/Y _16860_/X vssd1 vssd1 vccd1 vccd1 _25616_/A sky130_fd_sc_hd__a21oi_2
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18600_ _27689_/Q _18591_/X _18594_/X _18599_/Y vssd1 vssd1 vccd1 vccd1 _18600_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15812_ _13128_/X _26093_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15813_/A sky130_fd_sc_hd__mux2_1
X_19580_ _19580_/A vssd1 vssd1 vccd1 vccd1 _19580_/X sky130_fd_sc_hd__clkbuf_1
X_16792_ _16792_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _16793_/D sky130_fd_sc_hd__xnor2_1
XFILLER_19_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18531_ _26967_/Q _26935_/Q _26903_/Q _26871_/Q _18403_/X _18427_/X vssd1 vssd1 vccd1
+ vccd1 _18531_/X sky130_fd_sc_hd__mux4_1
X_15743_ _15743_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15743_/Y sky130_fd_sc_hd__nor2_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _15773_/A vssd1 vssd1 vccd1 vccd1 _13000_/A sky130_fd_sc_hd__clkbuf_2
X_27729_ _27729_/CLK _27729_/D vssd1 vssd1 vccd1 vccd1 _27729_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18462_ _18462_/A vssd1 vssd1 vccd1 vccd1 _18462_/X sky130_fd_sc_hd__buf_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _25655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15674_ _13184_/X _26147_/Q _15678_/S vssd1 vssd1 vccd1 vccd1 _15675_/A sky130_fd_sc_hd__mux2_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _27776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 _26819_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17413_ _17413_/A _17413_/B vssd1 vssd1 vccd1 vccd1 _17419_/A sky130_fd_sc_hd__or2_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14631_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_273 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_284 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18393_ _26544_/Q _26512_/Q _26480_/Q _27056_/Q _18392_/X _18259_/X vssd1 vssd1 vccd1
+ vccd1 _18393_/X sky130_fd_sc_hd__mux4_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17344_ _17299_/X _17337_/X _17340_/X _17343_/X vssd1 vssd1 vccd1 vccd1 _17344_/X
+ sky130_fd_sc_hd__o22a_1
X_14556_ _15716_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14556_/Y sky130_fd_sc_hd__nor2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13507_ _16495_/A vssd1 vssd1 vccd1 vccd1 _13900_/A sky130_fd_sc_hd__clkbuf_2
X_14487_ _15749_/A _14501_/B vssd1 vssd1 vccd1 vccd1 _14487_/Y sky130_fd_sc_hd__nor2_1
X_17275_ _17275_/A vssd1 vssd1 vccd1 vccd1 _27937_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19014_ _19113_/A _19014_/B vssd1 vssd1 vccd1 vccd1 _19014_/X sky130_fd_sc_hd__or2_1
X_13438_ _13859_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13438_/Y sky130_fd_sc_hd__nor2_1
X_16226_ _16180_/X _16221_/X _16223_/Y _16224_/X _16225_/X vssd1 vssd1 vccd1 vccd1
+ _16745_/A sky130_fd_sc_hd__o41a_1
XFILLER_173_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16157_ _16157_/A _16274_/B _16252_/C vssd1 vssd1 vccd1 vccd1 _16445_/A sky130_fd_sc_hd__and3_1
X_13369_ _14759_/A vssd1 vssd1 vccd1 vccd1 _13369_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15108_ _14798_/X _26398_/Q _15112_/S vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__mux2_1
X_16088_ _16077_/X _16602_/B _16087_/X vssd1 vssd1 vccd1 vccd1 _16088_/Y sky130_fd_sc_hd__a21oi_1
X_15039_ _26428_/Q _15028_/X _15029_/X _15038_/Y vssd1 vssd1 vccd1 vccd1 _26428_/D
+ sky130_fd_sc_hd__a31o_1
X_19916_ _25653_/A vssd1 vssd1 vccd1 vccd1 _20266_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19847_ _19847_/A vssd1 vssd1 vccd1 vccd1 _19847_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19778_ _19764_/X _19765_/X _19766_/X _19767_/X _19768_/X _19769_/X vssd1 vssd1 vccd1
+ vccd1 _19779_/A sky130_fd_sc_hd__mux4_1
XFILLER_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18729_ _26026_/Q _17728_/X _18735_/S vssd1 vssd1 vccd1 vccd1 _18730_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21740_ _21740_/A vssd1 vssd1 vccd1 vccd1 _21740_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21671_ _22543_/A vssd1 vssd1 vccd1 vccd1 _22019_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23410_ _23410_/A _23410_/B _23410_/C _23410_/D vssd1 vssd1 vccd1 vccd1 _23410_/Y
+ sky130_fd_sc_hd__nor4_1
X_20622_ _20708_/A vssd1 vssd1 vccd1 vccd1 _20687_/A sky130_fd_sc_hd__clkbuf_2
X_24390_ _24435_/A vssd1 vssd1 vccd1 vccd1 _24538_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23341_ _27767_/Q vssd1 vssd1 vccd1 vccd1 _24769_/A sky130_fd_sc_hd__clkinv_2
XFILLER_138_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20553_ _20601_/A vssd1 vssd1 vccd1 vccd1 _20553_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26060_ _26067_/CLK _26060_/D vssd1 vssd1 vccd1 vccd1 _26060_/Q sky130_fd_sc_hd__dfxtp_1
X_23272_ _27733_/Q vssd1 vssd1 vccd1 vccd1 _23272_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20484_ _20500_/A vssd1 vssd1 vccd1 vccd1 _20484_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25011_ _27231_/Q vssd1 vssd1 vccd1 vccd1 _25046_/S sky130_fd_sc_hd__buf_2
X_22223_ _22213_/X _22214_/X _22215_/X _22216_/X _22217_/X _22218_/X vssd1 vssd1 vccd1
+ vccd1 _22224_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22154_ _22154_/A vssd1 vssd1 vccd1 vccd1 _22154_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21105_ _21093_/X _21094_/X _21095_/X _21096_/X _21097_/X _21098_/X vssd1 vssd1 vccd1
+ vccd1 _21106_/A sky130_fd_sc_hd__mux4_1
X_22085_ _22085_/A vssd1 vssd1 vccd1 vccd1 _22085_/X sky130_fd_sc_hd__clkbuf_1
X_26962_ _22676_/X _26962_/D vssd1 vssd1 vccd1 vccd1 _26962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25913_ _25913_/CLK _25913_/D vssd1 vssd1 vccd1 vccd1 _25913_/Q sky130_fd_sc_hd__dfxtp_1
X_21036_ _21036_/A vssd1 vssd1 vccd1 vccd1 _21036_/X sky130_fd_sc_hd__clkbuf_1
X_26893_ _22430_/X _26893_/D vssd1 vssd1 vccd1 vccd1 _26893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25844_ _27130_/CLK _25844_/D vssd1 vssd1 vccd1 vccd1 _25844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25775_ _17479_/X _27843_/Q _25779_/S vssd1 vssd1 vccd1 vccd1 _25776_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22987_ _22974_/X _22976_/X _22978_/X _22980_/X _22981_/X _22982_/X vssd1 vssd1 vccd1
+ vccd1 _22988_/A sky130_fd_sc_hd__mux4_1
XFILLER_41_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27514_ _27515_/CLK _27514_/D vssd1 vssd1 vccd1 vccd1 _27514_/Q sky130_fd_sc_hd__dfxtp_1
X_21938_ _21986_/A vssd1 vssd1 vccd1 vccd1 _21938_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_24726_ _27607_/Q _24714_/X _24725_/X _24717_/X vssd1 vssd1 vccd1 vccd1 _27607_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24657_ _27581_/Q _24643_/X _24656_/X _24650_/X vssd1 vssd1 vccd1 vccd1 _27581_/D
+ sky130_fd_sc_hd__o211a_1
X_27445_ _27461_/CLK _27445_/D vssd1 vssd1 vccd1 vccd1 _27445_/Q sky130_fd_sc_hd__dfxtp_1
X_21869_ _21863_/X _21864_/X _21865_/X _21866_/X _21867_/X _21868_/X vssd1 vssd1 vccd1
+ vccd1 _21870_/A sky130_fd_sc_hd__mux4_1
XFILLER_179_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14410_/A _14412_/B vssd1 vssd1 vccd1 vccd1 _14410_/Y sky130_fd_sc_hd__nor2_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23608_ _24954_/B _27222_/Q _23616_/S vssd1 vssd1 vccd1 vccd1 _23609_/B sky130_fd_sc_hd__mux2_1
X_15390_ _14788_/X _26273_/Q _15390_/S vssd1 vssd1 vccd1 vccd1 _15391_/A sky130_fd_sc_hd__mux2_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24588_ _24588_/A vssd1 vssd1 vccd1 vccd1 _27554_/D sky130_fd_sc_hd__clkbuf_1
X_27376_ _27377_/CLK _27376_/D vssd1 vssd1 vccd1 vccd1 _27376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_772 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _26678_/Q _14337_/X _14329_/X _14340_/Y vssd1 vssd1 vccd1 vccd1 _26678_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23539_ _27761_/Q _27203_/Q _23542_/S vssd1 vssd1 vccd1 vccd1 _23540_/B sky130_fd_sc_hd__mux2_1
X_26327_ _20459_/X _26327_/D vssd1 vssd1 vccd1 vccd1 _26327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17060_ _17052_/X _17053_/X _17055_/X _17059_/X vssd1 vssd1 vccd1 vccd1 _17060_/X
+ sky130_fd_sc_hd__o22a_1
X_14272_ _14359_/A _14276_/B vssd1 vssd1 vccd1 vccd1 _14272_/Y sky130_fd_sc_hd__nor2_1
X_26258_ _20213_/X _26258_/D vssd1 vssd1 vccd1 vccd1 _26258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16011_ _27483_/Q _27270_/Q vssd1 vssd1 vccd1 vccd1 _16012_/B sky130_fd_sc_hd__xnor2_1
X_25209_ _27532_/Q _27500_/Q vssd1 vssd1 vccd1 vccd1 _25211_/A sky130_fd_sc_hd__nand2_1
X_13223_ _27037_/Q _13222_/X _13229_/S vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26189_ _19971_/X _26189_/D vssd1 vssd1 vccd1 vccd1 _26189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_533 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _27349_/Q _13061_/A _13081_/A _27317_/Q _13153_/X vssd1 vssd1 vccd1 vccd1
+ _16249_/A sky130_fd_sc_hd__a221o_1
XFILLER_3_841 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13085_/A vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__buf_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _26270_/Q _26238_/Q _26206_/Q _26174_/Q _17873_/X _17937_/X vssd1 vssd1 vccd1
+ vccd1 _17962_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19701_ _19701_/A vssd1 vssd1 vccd1 vccd1 _19701_/X sky130_fd_sc_hd__clkbuf_1
X_16913_ _16578_/Y _16913_/B vssd1 vssd1 vccd1 vccd1 _16915_/A sky130_fd_sc_hd__and2b_1
X_17893_ _17893_/A _17813_/X vssd1 vssd1 vccd1 vccd1 _17893_/X sky130_fd_sc_hd__or2b_1
Xrepeater408 _26048_/CLK vssd1 vssd1 vccd1 vccd1 _26047_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_77_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater419 _27392_/CLK vssd1 vssd1 vccd1 vccd1 _27394_/CLK sky130_fd_sc_hd__clkbuf_1
X_19632_ _19632_/A vssd1 vssd1 vccd1 vccd1 _19632_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16844_ _16844_/A _16844_/B _16844_/C _16844_/D vssd1 vssd1 vccd1 vccd1 _16844_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19563_ _26425_/Q _26393_/Q _26361_/Q _26329_/Q _18793_/X _18795_/X vssd1 vssd1 vccd1
+ vccd1 _19563_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16775_ _16734_/X _16733_/X _16785_/A _16774_/X vssd1 vssd1 vccd1 vccd1 _16776_/B
+ sky130_fd_sc_hd__o211ai_1
X_13987_ _14005_/A vssd1 vssd1 vccd1 vccd1 _13987_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18514_ _18512_/X _18513_/X _18514_/S vssd1 vssd1 vccd1 vccd1 _18514_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15726_ _26128_/Q _15721_/X _15713_/X _15725_/Y vssd1 vssd1 vccd1 vccd1 _26128_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1168 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _23650_/A vssd1 vssd1 vccd1 vccd1 _25075_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19494_ _19484_/X _19489_/X _19493_/X _19448_/X _19469_/X vssd1 vssd1 vccd1 vccd1
+ _19495_/C sky130_fd_sc_hd__a221o_1
XFILLER_179_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18445_ _18509_/A _18445_/B _18445_/C vssd1 vssd1 vccd1 vccd1 _18446_/A sky130_fd_sc_hd__and3_1
X_15657_ _15657_/A vssd1 vssd1 vccd1 vccd1 _26155_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _15769_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14608_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18376_ _27815_/Q _26576_/Q _26448_/Q _26128_/Q _18242_/X _18267_/X vssd1 vssd1 vccd1
+ vccd1 _18376_/X sky130_fd_sc_hd__mux4_2
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _26186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ input35/X vssd1 vssd1 vccd1 vccd1 _17370_/S sky130_fd_sc_hd__buf_2
XFILLER_186_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14539_ _26617_/Q _14530_/X _14536_/X _14538_/Y vssd1 vssd1 vccd1 vccd1 _26617_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _17238_/X _17253_/X _17255_/X _17257_/X vssd1 vssd1 vccd1 vccd1 _17258_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16209_ _26048_/Q _16221_/B _16221_/C vssd1 vssd1 vccd1 vccd1 _16209_/X sky130_fd_sc_hd__and3_1
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17189_ _27209_/Q _17188_/X _17189_/S vssd1 vssd1 vccd1 vccd1 _17190_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22910_ _22958_/A vssd1 vssd1 vccd1 vccd1 _22910_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23890_ _25926_/Q _25992_/Q _25825_/Q _26024_/Q _23852_/X _23882_/X vssd1 vssd1 vccd1
+ vccd1 _23890_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22841_ _22857_/A vssd1 vssd1 vccd1 vccd1 _22841_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25560_ _25560_/A vssd1 vssd1 vccd1 vccd1 _25560_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22772_ _22772_/A vssd1 vssd1 vccd1 vccd1 _22772_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24511_ _24511_/A vssd1 vssd1 vccd1 vccd1 _24589_/A sky130_fd_sc_hd__buf_2
X_21723_ _21739_/A vssd1 vssd1 vccd1 vccd1 _21723_/X sky130_fd_sc_hd__clkbuf_1
X_25491_ _27699_/Q _25479_/X _25480_/X vssd1 vssd1 vccd1 vccd1 _25491_/Y sky130_fd_sc_hd__a21oi_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27230_ _27826_/CLK _27230_/D vssd1 vssd1 vccd1 vccd1 _27230_/Q sky130_fd_sc_hd__dfxtp_1
X_24442_ _24442_/A vssd1 vssd1 vccd1 vccd1 _27498_/D sky130_fd_sc_hd__clkbuf_1
X_21654_ _21726_/A vssd1 vssd1 vccd1 vccd1 _21654_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27161_ _27420_/CLK _27161_/D vssd1 vssd1 vccd1 vccd1 _27161_/Q sky130_fd_sc_hd__dfxtp_1
X_20605_ _20673_/A vssd1 vssd1 vccd1 vccd1 _20605_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24373_ _24373_/A vssd1 vssd1 vccd1 vccd1 _27468_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21585_ _21585_/A vssd1 vssd1 vccd1 vccd1 _21650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26112_ _19705_/X _26112_/D vssd1 vssd1 vccd1 vccd1 _26112_/Q sky130_fd_sc_hd__dfxtp_1
X_23324_ input57/X input58/X input59/X input60/X vssd1 vssd1 vccd1 vccd1 _23325_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27092_ _27092_/CLK _27092_/D vssd1 vssd1 vccd1 vccd1 _27092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20536_ _20708_/A vssd1 vssd1 vccd1 vccd1 _20601_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26043_ _27356_/CLK _26043_/D vssd1 vssd1 vccd1 vccd1 _26043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23255_ _27737_/Q vssd1 vssd1 vccd1 vccd1 _23255_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_616 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20467_ _20515_/A vssd1 vssd1 vccd1 vccd1 _20467_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22206_ _22206_/A vssd1 vssd1 vccd1 vccd1 _22206_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23186_ _23186_/A vssd1 vssd1 vccd1 vccd1 _27130_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20398_ _20392_/X _20393_/X _20394_/X _20395_/X _20396_/X _20397_/X vssd1 vssd1 vccd1
+ vccd1 _20399_/A sky130_fd_sc_hd__mux4_1
XFILLER_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22137_ _22125_/X _22126_/X _22127_/X _22128_/X _22129_/X _22130_/X vssd1 vssd1 vccd1
+ vccd1 _22138_/A sky130_fd_sc_hd__mux4_1
XFILLER_160_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27994_ _27994_/A _15887_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
XFILLER_181_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22068_ _22084_/A vssd1 vssd1 vccd1 vccd1 _22068_/X sky130_fd_sc_hd__clkbuf_1
X_26945_ _22620_/X _26945_/D vssd1 vssd1 vccd1 vccd1 _26945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13910_ _13910_/A _13917_/B vssd1 vssd1 vccd1 vccd1 _13910_/Y sky130_fd_sc_hd__nor2_1
X_21019_ _21007_/X _21008_/X _21009_/X _21010_/X _21011_/X _21012_/X vssd1 vssd1 vccd1
+ vccd1 _21020_/A sky130_fd_sc_hd__mux4_1
XFILLER_87_472 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26876_ _22378_/X _26876_/D vssd1 vssd1 vccd1 vccd1 _26876_/Q sky130_fd_sc_hd__dfxtp_1
X_14890_ _14715_/X _26488_/Q _14896_/S vssd1 vssd1 vccd1 vccd1 _14891_/A sky130_fd_sc_hd__mux2_1
X_27987__453 vssd1 vssd1 vccd1 vccd1 _27987__453/HI _27987_/A sky130_fd_sc_hd__conb_1
X_13841_ _26845_/Q _13832_/X _13833_/X _13840_/Y vssd1 vssd1 vccd1 vccd1 _26845_/D
+ sky130_fd_sc_hd__a31o_1
X_25827_ _26026_/CLK _25827_/D vssd1 vssd1 vccd1 vccd1 _25827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13772_ _13779_/A vssd1 vssd1 vccd1 vccd1 _13827_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16560_ _16798_/A _16301_/B _16301_/C _16576_/A vssd1 vssd1 vccd1 vccd1 _16561_/B
+ sky130_fd_sc_hd__o31a_1
X_25758_ _25758_/A vssd1 vssd1 vccd1 vccd1 _27835_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15511_ _15511_/A vssd1 vssd1 vccd1 vccd1 _26220_/D sky130_fd_sc_hd__clkbuf_1
X_24709_ _27185_/Q _24711_/B vssd1 vssd1 vccd1 vccd1 _24709_/X sky130_fd_sc_hd__or2_1
XFILLER_71_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16491_ _16271_/A _16384_/X _16375_/B _25961_/Q _16490_/Y vssd1 vssd1 vccd1 vccd1
+ _16809_/B sky130_fd_sc_hd__a221o_2
XFILLER_167_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25689_ _25721_/A vssd1 vssd1 vccd1 vccd1 _25689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18230_ _18230_/A _18207_/X vssd1 vssd1 vccd1 vccd1 _18230_/X sky130_fd_sc_hd__or2b_1
X_27428_ _27437_/CLK _27428_/D vssd1 vssd1 vccd1 vccd1 _27428_/Q sky130_fd_sc_hd__dfxtp_1
X_15442_ _15464_/A vssd1 vssd1 vccd1 vccd1 _15451_/S sky130_fd_sc_hd__buf_2
XFILLER_169_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18161_ _18161_/A _18066_/X vssd1 vssd1 vccd1 vccd1 _18161_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15373_ _14763_/X _26281_/Q _15379_/S vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__mux2_1
X_27359_ _27478_/CLK _27359_/D vssd1 vssd1 vccd1 vccd1 _27359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17112_ _27074_/Q _27106_/Q _17112_/S vssd1 vssd1 vccd1 vccd1 _17112_/X sky130_fd_sc_hd__mux2_1
X_14324_ _26683_/Q _14322_/X _14248_/B _14323_/Y vssd1 vssd1 vccd1 vccd1 _26683_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18092_ _26147_/Q _26083_/Q _27011_/Q _26979_/Q _17821_/X _24386_/A vssd1 vssd1 vccd1
+ vccd1 _18093_/A sky130_fd_sc_hd__mux4_1
XFILLER_171_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14255_ _26709_/Q _14238_/X _14242_/X _14254_/Y vssd1 vssd1 vccd1 vccd1 _26709_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_116_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17043_ _17380_/S vssd1 vssd1 vccd1 vccd1 _17097_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _27040_/Q _13204_/X _13229_/S vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14186_ _14225_/A vssd1 vssd1 vccd1 vccd1 _14186_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13137_ _27352_/Q _13019_/A _13027_/A _27320_/Q _13136_/X vssd1 vssd1 vccd1 vccd1
+ _16271_/A sky130_fd_sc_hd__a221o_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18994_ _26816_/Q _26784_/Q _26752_/Q _26720_/Q _18870_/X _18967_/X vssd1 vssd1 vccd1
+ vccd1 _18995_/B sky130_fd_sc_hd__mux4_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17942_/X _17944_/X _18568_/S vssd1 vssd1 vccd1 vccd1 _17945_/X sky130_fd_sc_hd__mux2_1
X_13068_ _27063_/Q _13067_/X _13079_/S vssd1 vssd1 vccd1 vccd1 _13069_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater205 _25986_/CLK vssd1 vssd1 vccd1 vccd1 _25884_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater216 _27302_/CLK vssd1 vssd1 vccd1 vccd1 _27790_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_79_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater227 _26068_/CLK vssd1 vssd1 vccd1 vccd1 _25974_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater238 _27190_/CLK vssd1 vssd1 vccd1 vccd1 _27751_/CLK sky130_fd_sc_hd__clkbuf_1
X_17876_ _26523_/Q _26491_/Q _26459_/Q _27035_/Q _17841_/X _17843_/X vssd1 vssd1 vccd1
+ vccd1 _17876_/X sky130_fd_sc_hd__mux4_1
Xrepeater249 _27606_/CLK vssd1 vssd1 vccd1 vccd1 _27527_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19615_ _19605_/X _19606_/X _19607_/X _19608_/X _19609_/X _19610_/X vssd1 vssd1 vccd1
+ vccd1 _19616_/A sky130_fd_sc_hd__mux4_1
X_16827_ _16803_/Y _16825_/X _16826_/Y vssd1 vssd1 vccd1 vccd1 _16827_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19546_ _26552_/Q _26520_/Q _26488_/Q _27064_/Q _18896_/X _18898_/X vssd1 vssd1 vccd1
+ vccd1 _19546_/X sky130_fd_sc_hd__mux4_1
X_16758_ _16862_/A _16862_/B vssd1 vssd1 vccd1 vccd1 _16758_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_94_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15709_ _26134_/Q _15705_/X _15697_/X _15708_/Y vssd1 vssd1 vccd1 vccd1 _26134_/D
+ sky130_fd_sc_hd__a31o_1
X_19477_ _19431_/X _19476_/X _19387_/X vssd1 vssd1 vccd1 vccd1 _19477_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16689_ _16076_/A _16779_/A _16688_/Y _16699_/A vssd1 vssd1 vccd1 vccd1 _16689_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18428_ _26962_/Q _26930_/Q _26898_/Q _26866_/Q _18403_/X _18427_/X vssd1 vssd1 vccd1
+ vccd1 _18428_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18359_ _26831_/Q _26799_/Q _26767_/Q _26735_/Q _18358_/X _18199_/X vssd1 vssd1 vccd1
+ vccd1 _18359_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21370_ _21370_/A vssd1 vssd1 vccd1 vccd1 _21370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20321_ _20337_/A vssd1 vssd1 vccd1 vccd1 _20321_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23040_ _27066_/Q _17673_/X _23048_/S vssd1 vssd1 vccd1 vccd1 _23041_/A sky130_fd_sc_hd__mux2_1
X_20252_ _20338_/A vssd1 vssd1 vccd1 vccd1 _20322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20183_ _20249_/A vssd1 vssd1 vccd1 vccd1 _20183_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_547 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24991_ _25035_/A vssd1 vssd1 vccd1 vccd1 _24991_/X sky130_fd_sc_hd__buf_2
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26730_ _21870_/X _26730_/D vssd1 vssd1 vccd1 vccd1 _26730_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23942_ _23896_/X _23940_/X _23941_/X _23911_/X vssd1 vssd1 vccd1 vccd1 _27290_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26661_ _21624_/X _26661_/D vssd1 vssd1 vccd1 vccd1 _26661_/Q sky130_fd_sc_hd__dfxtp_1
X_23873_ _24014_/A vssd1 vssd1 vccd1 vccd1 _23873_/X sky130_fd_sc_hd__buf_2
XFILLER_45_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_25612_ _25547_/X _25552_/X _25553_/X _24970_/B _25554_/X vssd1 vssd1 vccd1 vccd1
+ _25612_/X sky130_fd_sc_hd__o311a_1
X_22824_ _22872_/A vssd1 vssd1 vccd1 vccd1 _22824_/X sky130_fd_sc_hd__clkbuf_1
X_26592_ _21384_/X _26592_/D vssd1 vssd1 vccd1 vccd1 _26592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25543_ _25543_/A vssd1 vssd1 vccd1 vccd1 _25543_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22755_ _22771_/A vssd1 vssd1 vccd1 vccd1 _22755_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21706_ _21738_/A vssd1 vssd1 vccd1 vccd1 _21706_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25474_ _25474_/A vssd1 vssd1 vccd1 vccd1 _25474_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22686_ _22686_/A vssd1 vssd1 vccd1 vccd1 _22686_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27213_ _27214_/CLK _27213_/D vssd1 vssd1 vccd1 vccd1 _27213_/Q sky130_fd_sc_hd__dfxtp_1
X_24425_ _27612_/Q _24433_/B vssd1 vssd1 vccd1 vccd1 _24426_/A sky130_fd_sc_hd__and2_1
X_21637_ _21631_/X _21632_/X _21633_/X _21634_/X _21635_/X _21636_/X vssd1 vssd1 vccd1
+ vccd1 _21638_/A sky130_fd_sc_hd__mux4_1
XFILLER_8_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27144_ _27144_/CLK _27144_/D vssd1 vssd1 vccd1 vccd1 _27144_/Q sky130_fd_sc_hd__dfxtp_1
X_24356_ _24356_/A vssd1 vssd1 vccd1 vccd1 _27460_/D sky130_fd_sc_hd__clkbuf_1
X_21568_ _21636_/A vssd1 vssd1 vccd1 vccd1 _21568_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23307_ _23306_/Y input53/X _23268_/Y input58/X vssd1 vssd1 vccd1 vccd1 _23307_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_20519_ _20587_/A vssd1 vssd1 vccd1 vccd1 _20519_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27075_ _27103_/CLK _27075_/D vssd1 vssd1 vccd1 vccd1 _27075_/Q sky130_fd_sc_hd__dfxtp_1
X_24287_ _24287_/A _24287_/B vssd1 vssd1 vccd1 vccd1 _24288_/A sky130_fd_sc_hd__and2_1
X_21499_ _21585_/A vssd1 vssd1 vccd1 vccd1 _21564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_154_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14040_ _14399_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14040_/Y sky130_fd_sc_hd__nor2_1
X_23238_ _23238_/A vssd1 vssd1 vccd1 vccd1 _27154_/D sky130_fd_sc_hd__clkbuf_1
X_26026_ _26026_/CLK _26026_/D vssd1 vssd1 vccd1 vccd1 _26026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23169_ _23169_/A vssd1 vssd1 vccd1 vccd1 _27123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27977_ _27977_/A _15908_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
X_15991_ _15991_/A vssd1 vssd1 vccd1 vccd1 _15992_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_612 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17730_ _17730_/A vssd1 vssd1 vccd1 vccd1 _25928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26928_ _22558_/X _26928_/D vssd1 vssd1 vccd1 vccd1 _26928_/Q sky130_fd_sc_hd__dfxtp_1
X_14942_ _14942_/A vssd1 vssd1 vccd1 vccd1 _14951_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17661_ _17508_/X _25901_/Q _17667_/S vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26859_ _22314_/X _26859_/D vssd1 vssd1 vccd1 vccd1 _26859_/Q sky130_fd_sc_hd__dfxtp_1
X_14873_ _26495_/Q _13405_/X _14879_/S vssd1 vssd1 vccd1 vccd1 _14874_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19400_ _26417_/Q _26385_/Q _26353_/Q _26321_/Q _19331_/X _19399_/X vssd1 vssd1 vccd1
+ vccd1 _19400_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16612_ _16077_/X _16783_/A _16611_/B _16087_/X vssd1 vssd1 vccd1 vccd1 _16612_/X
+ sky130_fd_sc_hd__a31o_1
X_13824_ _26852_/Q _13819_/X _13820_/X _13823_/Y vssd1 vssd1 vccd1 vccd1 _26852_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ _17592_/A vssd1 vssd1 vccd1 vccd1 _25870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19331_ _19465_/A vssd1 vssd1 vccd1 vccd1 _19331_/X sky130_fd_sc_hd__buf_2
X_16543_ _16494_/B _16500_/A _16494_/A vssd1 vssd1 vccd1 vccd1 _16543_/X sky130_fd_sc_hd__o21ba_1
XFILLER_16_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13755_ _13936_/A _13759_/B vssd1 vssd1 vccd1 vccd1 _13755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19262_ _26283_/Q _26251_/Q _26219_/Q _26187_/Q _19144_/X _19192_/X vssd1 vssd1 vccd1
+ vccd1 _19262_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16474_ _16772_/B vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13686_ _13740_/A vssd1 vssd1 vccd1 vccd1 _13698_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18213_ _26536_/Q _26504_/Q _26472_/Q _27048_/Q _18117_/X _18141_/X vssd1 vssd1 vccd1
+ vccd1 _18213_/X sky130_fd_sc_hd__mux4_1
X_15425_ _26258_/Q _13344_/X _15429_/S vssd1 vssd1 vccd1 vccd1 _15426_/A sky130_fd_sc_hd__mux2_1
X_19193_ _26280_/Q _26248_/Q _26216_/Q _26184_/Q _19144_/X _19192_/X vssd1 vssd1 vccd1
+ vccd1 _19193_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18144_ _18142_/X _18143_/X _18216_/S vssd1 vssd1 vccd1 vccd1 _18144_/X sky130_fd_sc_hd__mux2_1
X_15356_ _15356_/A vssd1 vssd1 vccd1 vccd1 _26289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_893 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14307_ _14396_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14307_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18075_ _18072_/X _18074_/X _18075_/S vssd1 vssd1 vccd1 vccd1 _18075_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15287_ _26319_/Q _13353_/X _15295_/S vssd1 vssd1 vccd1 vccd1 _15288_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17026_ _27196_/Q _17025_/X _17067_/S vssd1 vssd1 vccd1 vccd1 _17027_/A sky130_fd_sc_hd__mux2_1
X_14238_ _14296_/A vssd1 vssd1 vccd1 vccd1 _14238_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14169_ _26740_/Q _14157_/X _14167_/X _14168_/Y vssd1 vssd1 vccd1 vccd1 _26740_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18969_/X _18971_/X _18976_/X _18854_/X _18880_/X vssd1 vssd1 vccd1 vccd1
+ _18989_/B sky130_fd_sc_hd__a221o_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17928_ _18408_/A vssd1 vssd1 vccd1 vccd1 _17928_/X sky130_fd_sc_hd__clkbuf_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17859_ _17859_/A vssd1 vssd1 vccd1 vccd1 _25944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20870_ _20941_/A vssd1 vssd1 vccd1 vccd1 _20870_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19529_ _19527_/X _19528_/X _19565_/S vssd1 vssd1 vccd1 vccd1 _19529_/X sky130_fd_sc_hd__mux2_2
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22540_ _22540_/A vssd1 vssd1 vccd1 vccd1 _22889_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22471_ _22519_/A vssd1 vssd1 vccd1 vccd1 _22471_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24210_ _24210_/A _24210_/B vssd1 vssd1 vccd1 vccd1 _27374_/D sky130_fd_sc_hd__nor2_1
X_21422_ _21422_/A vssd1 vssd1 vccd1 vccd1 _21422_/X sky130_fd_sc_hd__clkbuf_1
X_25190_ _25190_/A _25190_/B vssd1 vssd1 vccd1 vccd1 _25191_/B sky130_fd_sc_hd__nand2_1
XFILLER_148_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24141_ _24141_/A vssd1 vssd1 vccd1 vccd1 _27343_/D sky130_fd_sc_hd__clkbuf_1
X_21353_ _21341_/X _21342_/X _21343_/X _21344_/X _21345_/X _21346_/X vssd1 vssd1 vccd1
+ vccd1 _21354_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20304_ _20336_/A vssd1 vssd1 vccd1 vccd1 _20304_/X sky130_fd_sc_hd__clkbuf_1
X_24072_ _27386_/Q _24072_/B vssd1 vssd1 vccd1 vccd1 _24073_/A sky130_fd_sc_hd__and2_1
X_21284_ _21284_/A vssd1 vssd1 vccd1 vccd1 _21284_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23023_ _23009_/X _23010_/X _23011_/X _23012_/X _23013_/X _23014_/X vssd1 vssd1 vccd1
+ vccd1 _23024_/A sky130_fd_sc_hd__mux4_1
XFILLER_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20235_ _20251_/A vssd1 vssd1 vccd1 vccd1 _20235_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27831_ _27832_/CLK _27831_/D vssd1 vssd1 vccd1 vccd1 _27831_/Q sky130_fd_sc_hd__dfxtp_1
X_20166_ _20338_/A vssd1 vssd1 vccd1 vccd1 _20236_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27762_ _27766_/CLK _27762_/D vssd1 vssd1 vccd1 vccd1 _27762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24974_ _27229_/Q vssd1 vssd1 vccd1 vccd1 _24974_/X sky130_fd_sc_hd__clkbuf_4
X_20097_ _20163_/A vssd1 vssd1 vccd1 vccd1 _20097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26713_ _21806_/X _26713_/D vssd1 vssd1 vccd1 vccd1 _26713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23925_ _23923_/X _23924_/X _23940_/S vssd1 vssd1 vccd1 vccd1 _23925_/X sky130_fd_sc_hd__mux2_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27693_ _27693_/CLK _27693_/D vssd1 vssd1 vccd1 vccd1 _27693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26644_ _21560_/X _26644_/D vssd1 vssd1 vccd1 vccd1 _26644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_648 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23856_ _24046_/S vssd1 vssd1 vccd1 vccd1 _23892_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22807_ _22893_/A vssd1 vssd1 vccd1 vccd1 _22872_/A sky130_fd_sc_hd__clkbuf_2
X_26575_ _21332_/X _26575_/D vssd1 vssd1 vccd1 vccd1 _26575_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_629 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20999_ _20991_/X _20992_/X _20993_/X _20994_/X _20995_/X _20996_/X vssd1 vssd1 vccd1
+ vccd1 _21000_/A sky130_fd_sc_hd__mux4_1
X_23787_ _25915_/Q _25981_/Q _25814_/Q _26013_/Q _23747_/X _23786_/X vssd1 vssd1 vccd1
+ vccd1 _23787_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25526_ _25500_/X _25230_/B _25525_/X _25513_/X vssd1 vssd1 vccd1 vccd1 _25526_/X
+ sky130_fd_sc_hd__a211o_1
X_13540_ _27344_/Q _13108_/X _13029_/A _27312_/Q _13182_/X vssd1 vssd1 vccd1 vccd1
+ _14500_/A sky130_fd_sc_hd__a221oi_4
XFILLER_164_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22738_ _22786_/A vssd1 vssd1 vccd1 vccd1 _22738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_201_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13878_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22669_ _22685_/A vssd1 vssd1 vccd1 vccd1 _22669_/X sky130_fd_sc_hd__clkbuf_2
X_25457_ _25456_/X _25440_/X _25442_/X _24838_/B _24384_/A vssd1 vssd1 vccd1 vccd1
+ _25457_/X sky130_fd_sc_hd__o311a_1
X_15210_ _14737_/X _26353_/Q _15212_/S vssd1 vssd1 vccd1 vccd1 _15211_/A sky130_fd_sc_hd__mux2_1
X_24408_ _24408_/A vssd1 vssd1 vccd1 vccd1 _27483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16190_ _23182_/B _16224_/B vssd1 vssd1 vccd1 vccd1 _16190_/Y sky130_fd_sc_hd__nor2_1
X_25388_ _25388_/A vssd1 vssd1 vccd1 vccd1 _27733_/D sky130_fd_sc_hd__clkbuf_1
X_27127_ _27127_/CLK _27127_/D vssd1 vssd1 vccd1 vccd1 _27127_/Q sky130_fd_sc_hd__dfxtp_1
X_15141_ _15141_/A vssd1 vssd1 vccd1 vccd1 _26384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24339_ _27553_/Q _24339_/B vssd1 vssd1 vccd1 vccd1 _24340_/A sky130_fd_sc_hd__and2_1
XFILLER_154_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15072_ _15072_/A vssd1 vssd1 vccd1 vccd1 _26415_/D sky130_fd_sc_hd__clkbuf_1
X_27058_ _23006_/X _27058_/D vssd1 vssd1 vccd1 vccd1 _27058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14023_ _14172_/A vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__clkbuf_2
X_18900_ _18922_/A vssd1 vssd1 vccd1 vccd1 _18900_/X sky130_fd_sc_hd__buf_6
X_26009_ _27109_/CLK _26009_/D vssd1 vssd1 vccd1 vccd1 _26009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19880_ _19866_/X _19867_/X _19868_/X _19869_/X _19870_/X _19871_/X vssd1 vssd1 vccd1
+ vccd1 _19881_/A sky130_fd_sc_hd__mux4_1
XFILLER_175_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18831_ _19287_/A vssd1 vssd1 vccd1 vccd1 _18831_/X sky130_fd_sc_hd__buf_2
XFILLER_68_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18762_ _18762_/A vssd1 vssd1 vccd1 vccd1 _26041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15974_ _15980_/A vssd1 vssd1 vccd1 vccd1 _15979_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17713_ _25923_/Q _17712_/X _17722_/S vssd1 vssd1 vccd1 vccd1 _17714_/A sky130_fd_sc_hd__mux2_1
X_14925_ _14766_/X _26472_/Q _14929_/S vssd1 vssd1 vccd1 vccd1 _14926_/A sky130_fd_sc_hd__mux2_1
X_18693_ _18761_/S vssd1 vssd1 vccd1 vccd1 _18702_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_49_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17644_ _17644_/A vssd1 vssd1 vccd1 vccd1 _25893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14856_ _14856_/A vssd1 vssd1 vccd1 vccd1 _26503_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13807_ _13833_/A vssd1 vssd1 vccd1 vccd1 _13807_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17575_ _17586_/A vssd1 vssd1 vccd1 vccd1 _17584_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14787_ _14787_/A vssd1 vssd1 vccd1 vccd1 _26530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19314_ _19314_/A vssd1 vssd1 vccd1 vccd1 _26061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16526_ _16908_/B _16526_/B vssd1 vssd1 vccd1 vccd1 _16552_/B sky130_fd_sc_hd__xor2_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13738_ _13917_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13738_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19245_ _19237_/X _19239_/X _19244_/X _19151_/X _19220_/X vssd1 vssd1 vccd1 vccd1
+ _19246_/C sky130_fd_sc_hd__a221o_2
XFILLER_176_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16457_ _27390_/Q _16457_/B vssd1 vssd1 vccd1 vccd1 _16457_/X sky130_fd_sc_hd__and2_1
X_13669_ _26907_/Q _13665_/X _13593_/B _13668_/Y vssd1 vssd1 vccd1 vccd1 _26907_/D
+ sky130_fd_sc_hd__a31o_1
X_15408_ _15464_/A vssd1 vssd1 vccd1 vccd1 _15477_/S sky130_fd_sc_hd__clkbuf_2
X_19176_ _19176_/A vssd1 vssd1 vccd1 vccd1 _26055_/D sky130_fd_sc_hd__clkbuf_1
X_16388_ _16388_/A vssd1 vssd1 vccd1 vccd1 _16747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18127_ _27804_/Q _26565_/Q _26437_/Q _26117_/Q _18099_/X _18126_/X vssd1 vssd1 vccd1
+ vccd1 _18127_/X sky130_fd_sc_hd__mux4_2
X_15339_ _15339_/A vssd1 vssd1 vccd1 vccd1 _26297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18058_ _18380_/A vssd1 vssd1 vccd1 vccd1 _18058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17009_ _23507_/A vssd1 vssd1 vccd1 vccd1 _25358_/B sky130_fd_sc_hd__buf_4
XFILLER_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20020_ _20009_/X _20011_/X _20013_/X _20015_/X _20016_/X _20017_/X vssd1 vssd1 vccd1
+ vccd1 _20021_/A sky130_fd_sc_hd__mux4_2
XFILLER_98_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1010 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21971_ _21965_/X _21966_/X _21967_/X _21968_/X _21969_/X _21970_/X vssd1 vssd1 vccd1
+ vccd1 _21972_/A sky130_fd_sc_hd__mux4_1
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23710_ _24947_/A _27259_/Q _23716_/S vssd1 vssd1 vccd1 vccd1 _23711_/A sky130_fd_sc_hd__mux2_1
X_20922_ _20954_/A vssd1 vssd1 vccd1 vccd1 _20922_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24690_ _24729_/A vssd1 vssd1 vccd1 vccd1 _24690_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23641_ _23641_/A vssd1 vssd1 vccd1 vccd1 _27230_/D sky130_fd_sc_hd__clkbuf_1
X_20853_ _20853_/A vssd1 vssd1 vccd1 vccd1 _20853_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23572_ _23572_/A vssd1 vssd1 vccd1 vccd1 _27212_/D sky130_fd_sc_hd__clkbuf_1
X_26360_ _20573_/X _26360_/D vssd1 vssd1 vccd1 vccd1 _26360_/Q sky130_fd_sc_hd__dfxtp_1
X_20784_ _20770_/X _20771_/X _20772_/X _20773_/X _20775_/X _20777_/X vssd1 vssd1 vccd1
+ vccd1 _20785_/A sky130_fd_sc_hd__mux4_1
XFILLER_195_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22523_ _22523_/A vssd1 vssd1 vccd1 vccd1 _22597_/A sky130_fd_sc_hd__buf_2
XFILLER_23_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25311_ _25329_/A _25329_/B _25304_/B vssd1 vssd1 vccd1 vccd1 _25312_/B sky130_fd_sc_hd__o21a_1
X_26291_ _20327_/X _26291_/D vssd1 vssd1 vccd1 vccd1 _26291_/Q sky130_fd_sc_hd__dfxtp_1
X_22454_ _22520_/A vssd1 vssd1 vccd1 vccd1 _22454_/X sky130_fd_sc_hd__clkbuf_1
X_25242_ _25266_/B _25242_/B vssd1 vssd1 vccd1 vccd1 _25243_/B sky130_fd_sc_hd__and2b_1
XFILLER_183_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21405_ _21389_/X _21390_/X _21391_/X _21392_/X _21394_/X _21396_/X vssd1 vssd1 vccd1
+ vccd1 _21406_/A sky130_fd_sc_hd__mux4_1
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25173_ _25173_/A _25173_/B vssd1 vssd1 vccd1 vccd1 _25174_/B sky130_fd_sc_hd__xnor2_1
XFILLER_109_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22385_ _22433_/A vssd1 vssd1 vccd1 vccd1 _22385_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24124_ _27441_/Q _24128_/B vssd1 vssd1 vccd1 vccd1 _24125_/A sky130_fd_sc_hd__and2_1
XFILLER_191_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21336_ _21336_/A vssd1 vssd1 vccd1 vccd1 _21336_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24055_ _25735_/B _24061_/B vssd1 vssd1 vccd1 vccd1 _24056_/A sky130_fd_sc_hd__and2_1
X_21267_ _21253_/X _21254_/X _21255_/X _21256_/X _21257_/X _21258_/X vssd1 vssd1 vccd1
+ vccd1 _21268_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23006_ _23006_/A vssd1 vssd1 vccd1 vccd1 _23006_/X sky130_fd_sc_hd__clkbuf_1
X_20218_ _20250_/A vssd1 vssd1 vccd1 vccd1 _20218_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21198_ _21214_/A vssd1 vssd1 vccd1 vccd1 _21198_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27814_ _25700_/X _27814_/D vssd1 vssd1 vccd1 vccd1 _27814_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ _20165_/A vssd1 vssd1 vccd1 vccd1 _20149_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_28012__478 vssd1 vssd1 vccd1 vccd1 _28012__478/HI _28012_/A sky130_fd_sc_hd__conb_1
XFILLER_92_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27745_ _27745_/CLK _27745_/D vssd1 vssd1 vccd1 vccd1 _27745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _12971_/A vssd1 vssd1 vccd1 vccd1 _27812_/D sky130_fd_sc_hd__clkbuf_1
X_24957_ _24962_/A _24957_/B vssd1 vssd1 vccd1 vccd1 _24957_/Y sky130_fd_sc_hd__nand2_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14710_ _14885_/A _15623_/B vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__or2_4
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23908_ _24002_/A vssd1 vssd1 vccd1 vccd1 _23908_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15690_ _15690_/A vssd1 vssd1 vccd1 vccd1 _26140_/D sky130_fd_sc_hd__clkbuf_1
X_27676_ _27676_/CLK _27676_/D vssd1 vssd1 vccd1 vccd1 _27967_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24888_ _24896_/C _24888_/B vssd1 vssd1 vccd1 vccd1 _24889_/B sky130_fd_sc_hd__or2_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26627_ _21508_/X _26627_/D vssd1 vssd1 vccd1 vccd1 _26627_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _15714_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23839_ _23837_/X _23838_/X _23846_/S vssd1 vssd1 vccd1 vccd1 _23839_/X sky130_fd_sc_hd__mux2_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17360_ _25941_/Q _26007_/Q _17370_/S vssd1 vssd1 vccd1 vccd1 _17361_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14572_ _26605_/Q _14563_/X _14566_/X _14571_/Y vssd1 vssd1 vccd1 vccd1 _26605_/D
+ sky130_fd_sc_hd__a31o_1
X_26558_ _21266_/X _26558_/D vssd1 vssd1 vccd1 vccd1 _26558_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16311_ _16412_/A vssd1 vssd1 vccd1 vccd1 _16311_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _26951_/Q _13510_/X _13505_/X _13522_/Y vssd1 vssd1 vccd1 vccd1 _26951_/D
+ sky130_fd_sc_hd__a31o_1
X_25509_ _25539_/A vssd1 vssd1 vccd1 vccd1 _25509_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17291_ _17291_/A vssd1 vssd1 vccd1 vccd1 _17341_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26489_ _21022_/X _26489_/D vssd1 vssd1 vccd1 vccd1 _26489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19030_ _18954_/X _19029_/X _18958_/X vssd1 vssd1 vccd1 vccd1 _19030_/X sky130_fd_sc_hd__o21a_1
XFILLER_202_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16242_ _24284_/A _27531_/Q _16242_/S vssd1 vssd1 vccd1 vccd1 _16728_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13454_ _13870_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13454_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13385_ _14775_/A vssd1 vssd1 vccd1 vccd1 _13385_/X sky130_fd_sc_hd__clkbuf_4
X_16173_ _26043_/Q _16201_/A _16194_/C vssd1 vssd1 vccd1 vccd1 _16173_/X sky130_fd_sc_hd__and3_1
XFILLER_12_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15124_ _15124_/A vssd1 vssd1 vccd1 vccd1 _26392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19932_ _19918_/X _19921_/X _19924_/X _19927_/X _19928_/X _19929_/X vssd1 vssd1 vccd1
+ vccd1 _19933_/A sky130_fd_sc_hd__mux4_1
X_15055_ _14721_/X _26422_/Q _15057_/S vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__mux2_1
X_14006_ _16451_/A vssd1 vssd1 vccd1 vccd1 _14374_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19863_ _19863_/A vssd1 vssd1 vccd1 vccd1 _19863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18814_ _18929_/A vssd1 vssd1 vccd1 vccd1 _18814_/X sky130_fd_sc_hd__clkbuf_2
X_19794_ _19780_/X _19781_/X _19782_/X _19783_/X _19784_/X _19785_/X vssd1 vssd1 vccd1
+ vccd1 _19795_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18745_ _18745_/A vssd1 vssd1 vccd1 vccd1 _26033_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15957_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15957_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14908_ _14908_/A vssd1 vssd1 vccd1 vccd1 _26480_/D sky130_fd_sc_hd__clkbuf_1
X_18676_ _18676_/A vssd1 vssd1 vccd1 vccd1 _18685_/S sky130_fd_sc_hd__buf_2
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _15894_/A vssd1 vssd1 vccd1 vccd1 _15893_/A sky130_fd_sc_hd__buf_6
X_17627_ _17627_/A vssd1 vssd1 vccd1 vccd1 _25885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14839_ _14839_/A vssd1 vssd1 vccd1 vccd1 _26511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17558_ _17463_/X _25855_/Q _17562_/S vssd1 vssd1 vccd1 vccd1 _17559_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _14753_/A _16501_/X _16311_/X _25962_/Q _16508_/Y vssd1 vssd1 vccd1 vccd1
+ _16666_/B sky130_fd_sc_hd__a221o_2
XFILLER_177_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17489_ _17505_/A vssd1 vssd1 vccd1 vccd1 _17502_/S sky130_fd_sc_hd__buf_2
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19228_ _26698_/Q _26666_/Q _26634_/Q _26602_/Q _19179_/X _19227_/X vssd1 vssd1 vccd1
+ vccd1 _19228_/X sky130_fd_sc_hd__mux4_2
XFILLER_20_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19159_ _26695_/Q _26663_/Q _26631_/Q _26599_/Q _19015_/X _19087_/X vssd1 vssd1 vccd1
+ vccd1 _19159_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22170_ _22170_/A vssd1 vssd1 vccd1 vccd1 _22170_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21121_ _21109_/X _21110_/X _21111_/X _21112_/X _21113_/X _21114_/X vssd1 vssd1 vccd1
+ vccd1 _21122_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21052_ _21052_/A vssd1 vssd1 vccd1 vccd1 _21052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20003_ _20003_/A vssd1 vssd1 vccd1 vccd1 _20003_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25860_ _26007_/CLK _25860_/D vssd1 vssd1 vccd1 vccd1 _25860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24811_ _24811_/A _24815_/B vssd1 vssd1 vccd1 vccd1 _24811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_507 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25791_ _25791_/A vssd1 vssd1 vccd1 vccd1 _27850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27530_ _27531_/CLK _27530_/D vssd1 vssd1 vccd1 vccd1 _27530_/Q sky130_fd_sc_hd__dfxtp_2
X_24742_ _24771_/A vssd1 vssd1 vccd1 vccd1 _24742_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21954_ _21986_/A vssd1 vssd1 vccd1 vccd1 _21954_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20905_ _20953_/A vssd1 vssd1 vccd1 vccd1 _20905_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27461_ _27461_/CLK _27461_/D vssd1 vssd1 vccd1 vccd1 _27461_/Q sky130_fd_sc_hd__dfxtp_1
X_21885_ _21879_/X _21880_/X _21881_/X _21882_/X _21883_/X _21884_/X vssd1 vssd1 vccd1
+ vccd1 _21886_/A sky130_fd_sc_hd__mux4_1
XFILLER_199_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24673_ _24700_/A vssd1 vssd1 vccd1 vccd1 _24673_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26412_ _20749_/X _26412_/D vssd1 vssd1 vccd1 vccd1 _26412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20836_ _20852_/A vssd1 vssd1 vccd1 vccd1 _20836_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23624_ _23624_/A _23624_/B vssd1 vssd1 vccd1 vccd1 _23625_/A sky130_fd_sc_hd__and2_1
X_27392_ _27392_/CLK _27392_/D vssd1 vssd1 vccd1 vccd1 _27392_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_910 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26343_ _20509_/X _26343_/D vssd1 vssd1 vccd1 vccd1 _26343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20767_ _20767_/A vssd1 vssd1 vccd1 vccd1 _20767_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23555_ _23555_/A vssd1 vssd1 vccd1 vccd1 _27207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22506_ _22522_/A vssd1 vssd1 vccd1 vccd1 _22506_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26274_ _20265_/X _26274_/D vssd1 vssd1 vccd1 vccd1 _26274_/Q sky130_fd_sc_hd__dfxtp_1
X_23486_ _27187_/Q _23495_/B vssd1 vssd1 vccd1 vccd1 _23486_/X sky130_fd_sc_hd__or2_1
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20698_ _20684_/X _20685_/X _20686_/X _20687_/X _20689_/X _20691_/X vssd1 vssd1 vccd1
+ vccd1 _20699_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_28013_ _28013_/A _15976_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_22437_ _22523_/A vssd1 vssd1 vccd1 vccd1 _22507_/A sky130_fd_sc_hd__buf_2
X_25225_ _25220_/A _25220_/B _25218_/A vssd1 vssd1 vccd1 vccd1 _25229_/A sky130_fd_sc_hd__o21ai_1
XFILLER_182_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ _27346_/Q _13019_/A _13027_/A _27314_/Q _13169_/X vssd1 vssd1 vccd1 vccd1
+ _16157_/A sky130_fd_sc_hd__a221o_1
X_22368_ _22434_/A vssd1 vssd1 vccd1 vccd1 _22368_/X sky130_fd_sc_hd__clkbuf_1
X_25156_ _25149_/A _25146_/X _25149_/B _25147_/A vssd1 vssd1 vccd1 vccd1 _25157_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21319_ _21301_/X _21302_/X _21303_/X _21304_/X _21307_/X _21310_/X vssd1 vssd1 vccd1
+ vccd1 _21320_/A sky130_fd_sc_hd__mux4_1
X_24107_ _24107_/A vssd1 vssd1 vccd1 vccd1 _27328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25087_ _25085_/X _25086_/X _25087_/S vssd1 vssd1 vccd1 vccd1 _25087_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22299_ _22347_/A vssd1 vssd1 vccd1 vccd1 _22299_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24038_ _24036_/X _24037_/X _24045_/S vssd1 vssd1 vccd1 vccd1 _24038_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_995 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16860_ _16752_/A _16754_/A _16859_/X vssd1 vssd1 vccd1 vccd1 _16860_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15811_ _15811_/A vssd1 vssd1 vccd1 vccd1 _26094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16791_ _16835_/A _16791_/B vssd1 vssd1 vccd1 vccd1 _16793_/C sky130_fd_sc_hd__xnor2_1
XFILLER_120_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25989_ _25989_/CLK _25989_/D vssd1 vssd1 vccd1 vccd1 _25989_/Q sky130_fd_sc_hd__dfxtp_1
X_18530_ _27822_/Q _26583_/Q _26455_/Q _26135_/Q _18401_/X _18425_/X vssd1 vssd1 vccd1
+ vccd1 _18530_/X sky130_fd_sc_hd__mux4_1
X_15742_ _26122_/Q _15734_/X _15740_/X _15741_/Y vssd1 vssd1 vccd1 vccd1 _26122_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27728_ _27752_/CLK _27728_/D vssd1 vssd1 vccd1 vccd1 _27728_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _23650_/A vssd1 vssd1 vccd1 vccd1 _15773_/A sky130_fd_sc_hd__buf_4
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _26547_/Q _26515_/Q _26483_/Q _27059_/Q _18392_/X _18418_/X vssd1 vssd1 vccd1
+ vccd1 _18461_/X sky130_fd_sc_hd__mux4_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27659_ _27659_/CLK _27659_/D vssd1 vssd1 vccd1 vccd1 _27659_/Q sky130_fd_sc_hd__dfxtp_1
X_15673_ _15673_/A vssd1 vssd1 vccd1 vccd1 _26148_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _24611_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 _25659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ _27407_/Q _27406_/Q _27405_/Q _27404_/Q vssd1 vssd1 vccd1 vccd1 _17413_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA_252 _27168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14707_/B vssd1 vssd1 vccd1 vccd1 _14624_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_263 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18392_/A vssd1 vssd1 vccd1 vccd1 _18392_/X sky130_fd_sc_hd__buf_2
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_741 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17343_ _17303_/X _17341_/X _17342_/X vssd1 vssd1 vccd1 vccd1 _17343_/X sky130_fd_sc_hd__a21bo_1
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14555_ _26612_/Q _14549_/X _14553_/X _14554_/Y vssd1 vssd1 vccd1 vccd1 _26612_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _27351_/Q _13062_/A _13082_/A _27319_/Q _13142_/X vssd1 vssd1 vccd1 vccd1
+ _16495_/A sky130_fd_sc_hd__a221oi_4
X_17274_ _27216_/Q _17273_/X _17311_/S vssd1 vssd1 vccd1 vccd1 _17275_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14501_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19013_ _26817_/Q _26785_/Q _26753_/Q _26721_/Q _18870_/X _18967_/X vssd1 vssd1 vccd1
+ vccd1 _19014_/B sky130_fd_sc_hd__mux4_1
X_16225_ _27524_/Q _16172_/X vssd1 vssd1 vccd1 vccd1 _16225_/X sky130_fd_sc_hd__or2b_1
X_13437_ _16099_/A vssd1 vssd1 vccd1 vccd1 _13859_/A sky130_fd_sc_hd__clkbuf_2
X_16156_ _16805_/A vssd1 vssd1 vccd1 vccd1 _16824_/A sky130_fd_sc_hd__clkbuf_2
X_13368_ _13368_/A vssd1 vssd1 vccd1 vccd1 _26987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _15107_/A vssd1 vssd1 vccd1 vccd1 _26399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16087_ _16650_/A vssd1 vssd1 vccd1 vccd1 _16087_/X sky130_fd_sc_hd__clkbuf_2
X_13299_ _13299_/A vssd1 vssd1 vccd1 vccd1 _27011_/D sky130_fd_sc_hd__clkbuf_1
X_15038_ _15777_/A _15043_/B vssd1 vssd1 vccd1 vccd1 _15038_/Y sky130_fd_sc_hd__nor2_1
X_19915_ _19915_/A vssd1 vssd1 vccd1 vccd1 _19915_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19846_ _19831_/X _19833_/X _19835_/X _19837_/X _19838_/X _19839_/X vssd1 vssd1 vccd1
+ vccd1 _19847_/A sky130_fd_sc_hd__mux4_1
XFILLER_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19777_ _19777_/A vssd1 vssd1 vccd1 vccd1 _19777_/X sky130_fd_sc_hd__clkbuf_1
X_16989_ _17252_/A vssd1 vssd1 vccd1 vccd1 _16989_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18728_ _18728_/A vssd1 vssd1 vccd1 vccd1 _26025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18659_ _25995_/Q _17731_/X _18663_/S vssd1 vssd1 vccd1 vccd1 _18660_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21670_ _21738_/A vssd1 vssd1 vccd1 vccd1 _21670_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20621_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20621_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23340_ _27769_/Q vssd1 vssd1 vccd1 vccd1 _24776_/A sky130_fd_sc_hd__clkinv_2
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20552_ _20600_/A vssd1 vssd1 vccd1 vccd1 _20552_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23271_ input67/X vssd1 vssd1 vccd1 vccd1 _23271_/Y sky130_fd_sc_hd__inv_2
X_20483_ _20515_/A vssd1 vssd1 vccd1 vccd1 _20483_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22222_ _22222_/A vssd1 vssd1 vccd1 vccd1 _22222_/X sky130_fd_sc_hd__clkbuf_1
X_25010_ _25916_/Q _25982_/Q _25815_/Q _26014_/Q _25009_/X _24983_/X vssd1 vssd1 vccd1
+ vccd1 _25010_/X sky130_fd_sc_hd__mux4_1
XFILLER_180_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22153_ _22141_/X _22142_/X _22143_/X _22144_/X _22145_/X _22146_/X vssd1 vssd1 vccd1
+ vccd1 _22154_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21104_ _21104_/A vssd1 vssd1 vccd1 vccd1 _21104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22084_ _22084_/A vssd1 vssd1 vccd1 vccd1 _22084_/X sky130_fd_sc_hd__clkbuf_1
X_26961_ _22674_/X _26961_/D vssd1 vssd1 vccd1 vccd1 _26961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_481 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25912_ _25913_/CLK _25912_/D vssd1 vssd1 vccd1 vccd1 _25912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21035_ _21023_/X _21024_/X _21025_/X _21026_/X _21027_/X _21028_/X vssd1 vssd1 vccd1
+ vccd1 _21036_/A sky130_fd_sc_hd__mux4_1
X_26892_ _22428_/X _26892_/D vssd1 vssd1 vccd1 vccd1 _26892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25843_ _27792_/CLK _25843_/D vssd1 vssd1 vccd1 vccd1 _25843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25774_ _25774_/A vssd1 vssd1 vccd1 vccd1 _27842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22986_ _22986_/A vssd1 vssd1 vccd1 vccd1 _22986_/X sky130_fd_sc_hd__clkbuf_1
X_27513_ _27515_/CLK _27513_/D vssd1 vssd1 vccd1 vccd1 _27513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24725_ _27191_/Q _24725_/B vssd1 vssd1 vccd1 vccd1 _24725_/X sky130_fd_sc_hd__or2_1
XFILLER_83_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21937_ _21985_/A vssd1 vssd1 vccd1 vccd1 _21937_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27444_ _27468_/CLK _27444_/D vssd1 vssd1 vccd1 vccd1 _27444_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24656_ _27165_/Q _24658_/B vssd1 vssd1 vccd1 vccd1 _24656_/X sky130_fd_sc_hd__or2_1
X_21868_ _21900_/A vssd1 vssd1 vccd1 vccd1 _21868_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23607_ _27780_/Q vssd1 vssd1 vccd1 vccd1 _24954_/B sky130_fd_sc_hd__buf_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27375_ _27787_/CLK _27375_/D vssd1 vssd1 vccd1 vccd1 _27375_/Q sky130_fd_sc_hd__dfxtp_1
X_20819_ _20867_/A vssd1 vssd1 vccd1 vccd1 _20819_/X sky130_fd_sc_hd__clkbuf_1
X_21799_ _21793_/X _21794_/X _21795_/X _21796_/X _21797_/X _21798_/X vssd1 vssd1 vccd1
+ vccd1 _21800_/A sky130_fd_sc_hd__mux4_1
X_24587_ _27654_/Q _24587_/B vssd1 vssd1 vccd1 vccd1 _24588_/A sky130_fd_sc_hd__and2_1
XFILLER_196_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14340_ _14340_/A _14350_/B vssd1 vssd1 vccd1 vccd1 _14340_/Y sky130_fd_sc_hd__nor2_1
X_26326_ _20457_/X _26326_/D vssd1 vssd1 vccd1 vccd1 _26326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23538_ _23538_/A vssd1 vssd1 vccd1 vccd1 _27202_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_784 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14271_ _14311_/A vssd1 vssd1 vccd1 vccd1 _14271_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26257_ _20211_/X _26257_/D vssd1 vssd1 vccd1 vccd1 _26257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_647 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23469_ _23482_/A vssd1 vssd1 vccd1 vccd1 _23469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16010_ _16264_/B vssd1 vssd1 vccd1 vccd1 _16297_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_1154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25208_ _25205_/A _25205_/B _25203_/A vssd1 vssd1 vccd1 vccd1 _25212_/A sky130_fd_sc_hd__o21ai_1
X_13222_ _14801_/A vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26188_ _19969_/X _26188_/D vssd1 vssd1 vccd1 vccd1 _26188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25139_ _25139_/A _25139_/B vssd1 vssd1 vccd1 vccd1 _25139_/Y sky130_fd_sc_hd__nand2_1
X_13153_ _27285_/Q _13176_/B vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__and2_1
XFILLER_98_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_853 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13084_ _27361_/Q _13063_/A _13082_/X _27329_/Q _13083_/X vssd1 vssd1 vccd1 vccd1
+ _13085_/A sky130_fd_sc_hd__a221o_1
XFILLER_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17961_ _17961_/A _17935_/X vssd1 vssd1 vccd1 vccd1 _17961_/X sky130_fd_sc_hd__or2b_1
XFILLER_124_589 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_28018__484 vssd1 vssd1 vccd1 vccd1 _28018__484/HI _28018_/A sky130_fd_sc_hd__conb_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16912_ _16647_/X _16908_/Y _16909_/Y _16911_/Y _16877_/X vssd1 vssd1 vccd1 vccd1
+ _24255_/A sky130_fd_sc_hd__o32a_1
X_19700_ _19694_/X _19695_/X _19696_/X _19697_/X _19698_/X _19699_/X vssd1 vssd1 vccd1
+ vccd1 _19701_/A sky130_fd_sc_hd__mux4_1
X_17892_ _26684_/Q _26652_/Q _26620_/Q _26588_/Q _17865_/X _17810_/X vssd1 vssd1 vccd1
+ vccd1 _17893_/A sky130_fd_sc_hd__mux4_1
Xrepeater409 _26048_/CLK vssd1 vssd1 vccd1 vccd1 _26049_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19631_ _19621_/X _19622_/X _19623_/X _19624_/X _19625_/X _19626_/X vssd1 vssd1 vccd1
+ vccd1 _19632_/A sky130_fd_sc_hd__mux4_1
X_16843_ _16843_/A _16843_/B _16758_/Y vssd1 vssd1 vccd1 vccd1 _16844_/D sky130_fd_sc_hd__or3b_1
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19562_ _19485_/X _19561_/X _19488_/X vssd1 vssd1 vccd1 vccd1 _19562_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16774_ _16774_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16774_/X sky130_fd_sc_hd__xor2_1
X_13986_ _26799_/Q _13969_/X _13983_/X _13985_/Y vssd1 vssd1 vccd1 vccd1 _26799_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18513_ _26966_/Q _26934_/Q _26902_/Q _26870_/Q _17903_/X _17904_/X vssd1 vssd1 vccd1
+ vccd1 _18513_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15725_ _15725_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15725_/Y sky130_fd_sc_hd__nor2_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12937_ _13244_/B vssd1 vssd1 vccd1 vccd1 _23650_/A sky130_fd_sc_hd__buf_2
X_19493_ _19490_/X _19491_/X _19565_/S vssd1 vssd1 vccd1 vccd1 _19493_/X sky130_fd_sc_hd__mux2_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18444_ _18436_/X _18439_/X _18442_/X _18443_/X _18372_/X vssd1 vssd1 vccd1 vccd1
+ _18445_/C sky130_fd_sc_hd__a221o_1
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15656_ _13139_/X _26155_/Q _15656_/S vssd1 vssd1 vccd1 vccd1 _15657_/A sky130_fd_sc_hd__mux2_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _26592_/Q _14602_/X _14605_/X _14606_/Y vssd1 vssd1 vccd1 vccd1 _26592_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18375_ _18375_/A vssd1 vssd1 vccd1 vccd1 _25965_/D sky130_fd_sc_hd__clkbuf_1
X_15587_ _26186_/Q _14759_/A _15595_/S vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__mux2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17326_ _27852_/Q _27156_/Q _25901_/Q _25869_/Q _17325_/X _17313_/X vssd1 vssd1 vccd1
+ vccd1 _17326_/X sky130_fd_sc_hd__mux4_1
XFILLER_193_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ _15699_/A _14542_/B vssd1 vssd1 vccd1 vccd1 _14538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17257_ _17242_/X _17256_/X _17220_/X vssd1 vssd1 vccd1 vccd1 _17257_/X sky130_fd_sc_hd__a21bo_1
X_14469_ _15736_/A _14483_/B vssd1 vssd1 vccd1 vccd1 _14469_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16208_ _16180_/X _16202_/X _16204_/Y _16206_/X _16207_/X vssd1 vssd1 vccd1 vccd1
+ _16378_/A sky130_fd_sc_hd__o41a_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17188_ _17184_/X _17186_/X _17235_/S vssd1 vssd1 vccd1 vccd1 _17188_/X sky130_fd_sc_hd__mux2_2
XFILLER_127_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16139_ _27403_/Q _16144_/B _16138_/Y _13077_/A vssd1 vssd1 vccd1 vccd1 _16139_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_429 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1093 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19829_ _19829_/A vssd1 vssd1 vccd1 vccd1 _19829_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22840_ _22872_/A vssd1 vssd1 vccd1 vccd1 _22840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22771_ _22771_/A vssd1 vssd1 vccd1 vccd1 _22771_/X sky130_fd_sc_hd__clkbuf_2
X_24510_ _24510_/A vssd1 vssd1 vccd1 vccd1 _27525_/D sky130_fd_sc_hd__clkbuf_1
X_21722_ _21738_/A vssd1 vssd1 vccd1 vccd1 _21722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25490_ _24756_/A _25474_/X _25486_/Y _25489_/X _25467_/X vssd1 vssd1 vccd1 vccd1
+ _27762_/D sky130_fd_sc_hd__a221oi_1
XFILLER_80_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21653_ _21653_/A vssd1 vssd1 vccd1 vccd1 _21726_/A sky130_fd_sc_hd__clkbuf_2
X_24441_ _27619_/Q _24445_/B vssd1 vssd1 vccd1 vccd1 _24442_/A sky130_fd_sc_hd__and2_1
XFILLER_33_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27160_ _27160_/CLK _27160_/D vssd1 vssd1 vccd1 vccd1 _27160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20604_ _20776_/A vssd1 vssd1 vccd1 vccd1 _20673_/A sky130_fd_sc_hd__clkbuf_2
X_21584_ _21649_/A vssd1 vssd1 vccd1 vccd1 _21584_/X sky130_fd_sc_hd__clkbuf_1
X_24372_ _27568_/Q _24372_/B vssd1 vssd1 vccd1 vccd1 _24373_/A sky130_fd_sc_hd__and2_1
XFILLER_32_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26111_ _19703_/X _26111_/D vssd1 vssd1 vccd1 vccd1 _26111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23323_ input61/X input62/X input64/X input65/X vssd1 vssd1 vccd1 vccd1 _23325_/B
+ sky130_fd_sc_hd__or4_1
X_20535_ _20600_/A vssd1 vssd1 vccd1 vccd1 _20535_/X sky130_fd_sc_hd__clkbuf_1
X_27091_ _27124_/CLK _27091_/D vssd1 vssd1 vccd1 vccd1 _27091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26042_ _27328_/CLK _26042_/D vssd1 vssd1 vccd1 vccd1 _26042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23254_ _27727_/Q vssd1 vssd1 vccd1 vccd1 _23254_/Y sky130_fd_sc_hd__inv_2
X_20466_ _20514_/A vssd1 vssd1 vccd1 vccd1 _20466_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_628 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22205_ _22194_/X _22196_/X _22198_/X _22200_/X _22201_/X _22202_/X vssd1 vssd1 vccd1
+ vccd1 _22206_/A sky130_fd_sc_hd__mux4_1
X_23185_ _17408_/X _27130_/Q _23193_/S vssd1 vssd1 vccd1 vccd1 _23186_/A sky130_fd_sc_hd__mux2_1
X_20397_ _20413_/A vssd1 vssd1 vccd1 vccd1 _20397_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22136_ _22136_/A vssd1 vssd1 vccd1 vccd1 _22136_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27993_ _27993_/A _15889_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22067_ _22083_/A vssd1 vssd1 vccd1 vccd1 _22067_/X sky130_fd_sc_hd__clkbuf_1
X_26944_ _22608_/X _26944_/D vssd1 vssd1 vccd1 vccd1 _26944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21018_ _21018_/A vssd1 vssd1 vccd1 vccd1 _21018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26875_ _22376_/X _26875_/D vssd1 vssd1 vccd1 vccd1 _26875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_484 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13840_ _13934_/A _13847_/B vssd1 vssd1 vccd1 vccd1 _13840_/Y sky130_fd_sc_hd__nor2_1
X_25826_ _27083_/CLK _25826_/D vssd1 vssd1 vccd1 vccd1 _25826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13771_ _26871_/Q _13761_/X _13764_/X _13770_/Y vssd1 vssd1 vccd1 vccd1 _26871_/D
+ sky130_fd_sc_hd__a31o_1
X_25757_ _17453_/X _27835_/Q _25757_/S vssd1 vssd1 vccd1 vccd1 _25758_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22969_ _22955_/X _22956_/X _22957_/X _22958_/X _22960_/X _22962_/X vssd1 vssd1 vccd1
+ vccd1 _22970_/A sky130_fd_sc_hd__mux4_1
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15510_ _13133_/X _26220_/Q _15512_/S vssd1 vssd1 vccd1 vccd1 _15511_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24708_ _24403_/A _24700_/X _24707_/X _24703_/X vssd1 vssd1 vccd1 vccd1 _27600_/D
+ sky130_fd_sc_hd__o211a_1
X_16490_ _16490_/A _16490_/B vssd1 vssd1 vccd1 vccd1 _16490_/Y sky130_fd_sc_hd__nor2_1
X_25688_ _25688_/A vssd1 vssd1 vccd1 vccd1 _25688_/X sky130_fd_sc_hd__clkbuf_1
X_27427_ _27427_/CLK _27427_/D vssd1 vssd1 vccd1 vccd1 _27427_/Q sky130_fd_sc_hd__dfxtp_1
X_15441_ _15441_/A vssd1 vssd1 vccd1 vccd1 _26251_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24639_ _24639_/A vssd1 vssd1 vccd1 vccd1 _27577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18160_ _26150_/Q _26086_/Q _27014_/Q _26982_/Q _18041_/X _18112_/X vssd1 vssd1 vccd1
+ vccd1 _18161_/A sky130_fd_sc_hd__mux4_1
X_15372_ _15372_/A vssd1 vssd1 vccd1 vccd1 _26282_/D sky130_fd_sc_hd__clkbuf_1
X_27358_ _27358_/CLK _27358_/D vssd1 vssd1 vccd1 vccd1 _27358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17111_ _17052_/X _17105_/X _17107_/X _17110_/X vssd1 vssd1 vccd1 vccd1 _17111_/X
+ sky130_fd_sc_hd__o22a_1
X_14323_ _14410_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14323_/Y sky130_fd_sc_hd__nor2_1
X_26309_ _20391_/X _26309_/D vssd1 vssd1 vccd1 vccd1 _26309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18091_ _18089_/X _18090_/X _18522_/S vssd1 vssd1 vccd1 vccd1 _18091_/X sky130_fd_sc_hd__mux2_1
X_27289_ _27423_/CLK _27289_/D vssd1 vssd1 vccd1 vccd1 _27289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17042_ _17029_/X _17042_/B vssd1 vssd1 vccd1 vccd1 _17042_/X sky130_fd_sc_hd__and2b_1
X_14254_ _14342_/A _14263_/B vssd1 vssd1 vccd1 vccd1 _14254_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_466 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13205_ _13205_/A vssd1 vssd1 vccd1 vccd1 _13229_/S sky130_fd_sc_hd__clkbuf_2
X_14185_ _26734_/Q _14173_/X _14181_/X _14184_/Y vssd1 vssd1 vccd1 vccd1 _26734_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13136_ _27288_/Q _13169_/B vssd1 vssd1 vccd1 vccd1 _13136_/X sky130_fd_sc_hd__and2_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18993_ _19428_/A vssd1 vssd1 vccd1 vccd1 _19113_/A sky130_fd_sc_hd__clkbuf_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _26397_/Q _26365_/Q _26333_/Q _26301_/Q _17877_/X _17943_/X vssd1 vssd1 vccd1
+ vccd1 _17944_/X sky130_fd_sc_hd__mux4_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13067_ _14718_/A vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__buf_2
XFILLER_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater206 _25987_/CLK vssd1 vssd1 vccd1 vccd1 _27140_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater217 _27302_/CLK vssd1 vssd1 vccd1 vccd1 _27789_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater228 _26067_/CLK vssd1 vssd1 vccd1 vccd1 _26068_/CLK sky130_fd_sc_hd__clkbuf_1
X_17875_ _17830_/X _17874_/X _17838_/X vssd1 vssd1 vccd1 vccd1 _17875_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater239 _27607_/CLK vssd1 vssd1 vccd1 vccd1 _27190_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19614_ _19614_/A vssd1 vssd1 vccd1 vccd1 _19614_/X sky130_fd_sc_hd__clkbuf_1
X_16826_ _16826_/A _16908_/B vssd1 vssd1 vccd1 vccd1 _16826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16757_ _16755_/Y _16756_/X _16753_/A vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__a21o_1
X_19545_ _26424_/Q _26392_/Q _26360_/Q _26328_/Q _19465_/X _18795_/X vssd1 vssd1 vccd1
+ vccd1 _19545_/X sky130_fd_sc_hd__mux4_1
X_13969_ _14005_/A vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_595 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15708_ _15708_/A _15718_/B vssd1 vssd1 vccd1 vccd1 _15708_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19476_ _26709_/Q _26677_/Q _26645_/Q _26613_/Q _18816_/X _19385_/X vssd1 vssd1 vccd1
+ vccd1 _19476_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16688_ _16779_/B vssd1 vssd1 vccd1 vccd1 _16688_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _18427_/A vssd1 vssd1 vccd1 vccd1 _18427_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15639_ _13094_/X _26163_/Q _15645_/S vssd1 vssd1 vccd1 vccd1 _15640_/A sky130_fd_sc_hd__mux2_1
X_18358_ _18358_/A vssd1 vssd1 vccd1 vccd1 _18358_/X sky130_fd_sc_hd__buf_2
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17309_ input38/X vssd1 vssd1 vccd1 vccd1 _17356_/S sky130_fd_sc_hd__clkbuf_2
X_18289_ _27811_/Q _26572_/Q _26444_/Q _26124_/Q _17996_/X _17997_/X vssd1 vssd1 vccd1
+ vccd1 _18289_/X sky130_fd_sc_hd__mux4_2
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20320_ _20336_/A vssd1 vssd1 vccd1 vccd1 _20320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20251_ _20251_/A vssd1 vssd1 vccd1 vccd1 _20251_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20182_ _20268_/A vssd1 vssd1 vccd1 vccd1 _20249_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24990_ _24990_/A vssd1 vssd1 vccd1 vccd1 _27673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23941_ _27085_/Q _23907_/X _23908_/X _27117_/Q _23909_/X vssd1 vssd1 vccd1 vccd1
+ _23941_/X sky130_fd_sc_hd__a221o_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26660_ _21622_/X _26660_/D vssd1 vssd1 vccd1 vccd1 _26660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23872_ _23849_/X _23870_/X _23871_/X _23864_/X vssd1 vssd1 vccd1 vccd1 _27282_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_454 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25611_ _27720_/Q _25539_/X _25540_/X vssd1 vssd1 vccd1 vccd1 _25611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22823_ _22871_/A vssd1 vssd1 vccd1 vccd1 _22823_/X sky130_fd_sc_hd__clkbuf_1
X_26591_ _21382_/X _26591_/D vssd1 vssd1 vccd1 vccd1 _26591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25542_ _25517_/X _25522_/X _25523_/X _24907_/B _25524_/X vssd1 vssd1 vccd1 vccd1
+ _25542_/X sky130_fd_sc_hd__o311a_1
XFILLER_53_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22754_ _22786_/A vssd1 vssd1 vccd1 vccd1 _22754_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21705_ _21737_/A vssd1 vssd1 vccd1 vccd1 _21705_/X sky130_fd_sc_hd__clkbuf_1
X_25473_ _24750_/A _25431_/X _25469_/Y _25472_/X _25467_/X vssd1 vssd1 vccd1 vccd1
+ _27759_/D sky130_fd_sc_hd__a221oi_1
X_22685_ _22685_/A vssd1 vssd1 vccd1 vccd1 _22685_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27212_ _27856_/CLK _27212_/D vssd1 vssd1 vccd1 vccd1 _27212_/Q sky130_fd_sc_hd__dfxtp_1
X_24424_ _24538_/A vssd1 vssd1 vccd1 vccd1 _24433_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21636_ _21636_/A vssd1 vssd1 vccd1 vccd1 _21636_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27143_ _27840_/CLK _27143_/D vssd1 vssd1 vccd1 vccd1 _27143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24355_ _27560_/Q _24361_/B vssd1 vssd1 vccd1 vccd1 _24356_/A sky130_fd_sc_hd__and2_1
XFILLER_193_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21567_ _21653_/A vssd1 vssd1 vccd1 vccd1 _21636_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23306_ _27741_/Q vssd1 vssd1 vccd1 vccd1 _23306_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20518_ _20776_/A vssd1 vssd1 vccd1 vccd1 _20587_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_27074_ _27135_/CLK _27074_/D vssd1 vssd1 vccd1 vccd1 _27074_/Q sky130_fd_sc_hd__dfxtp_1
X_21498_ _21563_/A vssd1 vssd1 vccd1 vccd1 _21498_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24286_ _16243_/Y _16244_/X _16245_/X _24279_/X vssd1 vssd1 vccd1 vccd1 _27421_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_119_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26025_ _27115_/CLK _26025_/D vssd1 vssd1 vccd1 vccd1 _26025_/Q sky130_fd_sc_hd__dfxtp_1
X_23237_ _17501_/X _27154_/Q _23237_/S vssd1 vssd1 vccd1 vccd1 _23238_/A sky130_fd_sc_hd__mux2_1
X_20449_ _20514_/A vssd1 vssd1 vccd1 vccd1 _20449_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23168_ _27123_/Q _17756_/X _23176_/S vssd1 vssd1 vccd1 vccd1 _23169_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22119_ _22103_/X _22106_/X _22109_/X _22112_/X _22113_/X _22114_/X vssd1 vssd1 vccd1
+ vccd1 _22120_/A sky130_fd_sc_hd__mux4_1
X_23099_ _27093_/Q _17763_/X _23103_/S vssd1 vssd1 vccd1 vccd1 _23100_/A sky130_fd_sc_hd__mux2_1
X_27976_ _27976_/A _15909_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_15990_ _27576_/Q vssd1 vssd1 vccd1 vccd1 _15991_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26927_ _22556_/X _26927_/D vssd1 vssd1 vccd1 vccd1 _26927_/Q sky130_fd_sc_hd__dfxtp_1
X_14941_ _14941_/A vssd1 vssd1 vccd1 vccd1 _26465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17660_ _17660_/A vssd1 vssd1 vccd1 vccd1 _25900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26858_ _22312_/X _26858_/D vssd1 vssd1 vccd1 vccd1 _26858_/Q sky130_fd_sc_hd__dfxtp_1
X_14872_ _14872_/A vssd1 vssd1 vccd1 vccd1 _26496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16611_ _16783_/A _16611_/B vssd1 vssd1 vccd1 vccd1 _16611_/X sky130_fd_sc_hd__or2_1
X_13823_ _13915_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13823_/Y sky130_fd_sc_hd__nor2_1
X_25809_ _25721_/X _25722_/X _25723_/X _25724_/X _25725_/X _25726_/X vssd1 vssd1 vccd1
+ vccd1 _25810_/A sky130_fd_sc_hd__mux4_2
X_17591_ _17511_/X _25870_/Q _17595_/S vssd1 vssd1 vccd1 vccd1 _17592_/A sky130_fd_sc_hd__mux2_1
X_26789_ _22066_/X _26789_/D vssd1 vssd1 vccd1 vccd1 _26789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ _16662_/A _16911_/A _16660_/A _16885_/A vssd1 vssd1 vccd1 vccd1 _16542_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19330_ _19191_/X _19329_/X _19194_/X vssd1 vssd1 vccd1 vccd1 _19330_/X sky130_fd_sc_hd__o21a_1
X_13754_ _26877_/Q _13750_/X _13745_/X _13753_/Y vssd1 vssd1 vccd1 vccd1 _26877_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_71_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19261_ _19261_/A _19261_/B vssd1 vssd1 vccd1 vccd1 _19261_/X sky130_fd_sc_hd__or2_1
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16473_ _16692_/B _16610_/A _16692_/C _16469_/X _16472_/X vssd1 vssd1 vccd1 vccd1
+ _16482_/B sky130_fd_sc_hd__a311o_1
X_13685_ _13691_/A vssd1 vssd1 vccd1 vccd1 _13740_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18212_ _18162_/X _18210_/X _18211_/X vssd1 vssd1 vccd1 vccd1 _18212_/X sky130_fd_sc_hd__o21a_1
X_15424_ _15424_/A vssd1 vssd1 vccd1 vccd1 _26259_/D sky130_fd_sc_hd__clkbuf_1
X_19192_ _19385_/A vssd1 vssd1 vccd1 vccd1 _19192_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18143_ _26405_/Q _26373_/Q _26341_/Q _26309_/Q _18048_/X _18073_/X vssd1 vssd1 vccd1
+ vccd1 _18143_/X sky130_fd_sc_hd__mux4_1
XFILLER_54_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15355_ _14737_/X _26289_/Q _15357_/S vssd1 vssd1 vccd1 vccd1 _15356_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ _26690_/Q _14296_/X _14297_/X _14305_/Y vssd1 vssd1 vccd1 vccd1 _26690_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18074_ _26402_/Q _26370_/Q _26338_/Q _26306_/Q _18048_/X _18073_/X vssd1 vssd1 vccd1
+ vccd1 _18074_/X sky130_fd_sc_hd__mux4_1
XFILLER_116_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15286_ _15332_/S vssd1 vssd1 vccd1 vccd1 _15295_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17025_ _17023_/X _17024_/X _17048_/S vssd1 vssd1 vccd1 vccd1 _17025_/X sky130_fd_sc_hd__mux2_1
X_14237_ _14548_/A vssd1 vssd1 vccd1 vccd1 _14296_/A sky130_fd_sc_hd__clkbuf_2
X_14168_ _14346_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_981 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13119_/A vssd1 vssd1 vccd1 vccd1 _27055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_557 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _26765_/Q _14090_/X _14093_/X _14098_/Y vssd1 vssd1 vccd1 vccd1 _26765_/D
+ sky130_fd_sc_hd__a31o_1
X_18976_ _18973_/X _18975_/X _19047_/S vssd1 vssd1 vccd1 vccd1 _18976_/X sky130_fd_sc_hd__mux2_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _26813_/Q _26781_/Q _26749_/Q _26717_/Q _17863_/X _17890_/X vssd1 vssd1 vccd1
+ vccd1 _17927_/X sky130_fd_sc_hd__mux4_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17858_ _24624_/B _17858_/B _17858_/C vssd1 vssd1 vccd1 vccd1 _17859_/A sky130_fd_sc_hd__and3_1
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16809_ _16809_/A _16809_/B vssd1 vssd1 vccd1 vccd1 _16809_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17789_ _18401_/A vssd1 vssd1 vccd1 vccd1 _17789_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_198_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19528_ _26551_/Q _26519_/Q _26487_/Q _27063_/Q _18896_/X _19445_/X vssd1 vssd1 vccd1
+ vccd1 _19528_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19459_ _19453_/X _19455_/X _19458_/X _18837_/X _19393_/X vssd1 vssd1 vccd1 vccd1
+ _19471_/B sky130_fd_sc_hd__a221o_1
XFILLER_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22470_ _22470_/A vssd1 vssd1 vccd1 vccd1 _22470_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21421_ _21408_/X _21410_/X _21412_/X _21414_/X _21415_/X _21416_/X vssd1 vssd1 vccd1
+ vccd1 _21422_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21352_ _21352_/A vssd1 vssd1 vccd1 vccd1 _21352_/X sky130_fd_sc_hd__clkbuf_1
X_24140_ _27448_/Q _24140_/B vssd1 vssd1 vccd1 vccd1 _24141_/A sky130_fd_sc_hd__and2_1
XFILLER_190_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20303_ _20335_/A vssd1 vssd1 vccd1 vccd1 _20303_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21283_ _21269_/X _21270_/X _21271_/X _21272_/X _21273_/X _21274_/X vssd1 vssd1 vccd1
+ vccd1 _21284_/A sky130_fd_sc_hd__mux4_1
X_24071_ _24071_/A vssd1 vssd1 vccd1 vccd1 _27312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20234_ _20250_/A vssd1 vssd1 vccd1 vccd1 _20234_/X sky130_fd_sc_hd__clkbuf_1
X_23022_ _23022_/A vssd1 vssd1 vccd1 vccd1 _23022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27830_ _27830_/CLK _27830_/D vssd1 vssd1 vccd1 vccd1 _27830_/Q sky130_fd_sc_hd__dfxtp_1
X_20165_ _20165_/A vssd1 vssd1 vccd1 vccd1 _20165_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_27761_ _27766_/CLK _27761_/D vssd1 vssd1 vccd1 vccd1 _27761_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24973_ _27826_/Q _27130_/Q _25875_/Q _25843_/Q _24972_/X _23638_/B vssd1 vssd1 vccd1
+ vccd1 _24973_/X sky130_fd_sc_hd__mux4_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20096_ _20268_/A vssd1 vssd1 vccd1 vccd1 _20163_/A sky130_fd_sc_hd__buf_2
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26712_ _21804_/X _26712_/D vssd1 vssd1 vccd1 vccd1 _26712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23924_ _27083_/Q _27115_/Q _23939_/S vssd1 vssd1 vccd1 vccd1 _23924_/X sky130_fd_sc_hd__mux2_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27692_ _27695_/CLK _27692_/D vssd1 vssd1 vccd1 vccd1 _27692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26643_ _21558_/X _26643_/D vssd1 vssd1 vccd1 vccd1 _26643_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23855_ _23851_/X _23853_/X _23891_/S vssd1 vssd1 vccd1 vccd1 _23855_/X sky130_fd_sc_hd__mux2_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22806_ _22871_/A vssd1 vssd1 vccd1 vccd1 _22806_/X sky130_fd_sc_hd__clkbuf_1
X_26574_ _21320_/X _26574_/D vssd1 vssd1 vccd1 vccd1 _26574_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23786_ _23929_/A vssd1 vssd1 vccd1 vccd1 _23786_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20998_ _20998_/A vssd1 vssd1 vccd1 vccd1 _20998_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25525_ _25517_/X _25522_/X _25523_/X _24894_/B _25524_/X vssd1 vssd1 vccd1 vccd1
+ _25525_/X sky130_fd_sc_hd__o311a_1
XFILLER_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22737_ _22785_/A vssd1 vssd1 vccd1 vccd1 _22737_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _16563_/A vssd1 vssd1 vccd1 vccd1 _13878_/A sky130_fd_sc_hd__clkbuf_2
X_25456_ _25517_/A vssd1 vssd1 vccd1 vccd1 _25456_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22668_ _22700_/A vssd1 vssd1 vccd1 vccd1 _22668_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_528 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24407_ _24407_/A _24411_/B vssd1 vssd1 vccd1 vccd1 _24408_/A sky130_fd_sc_hd__and2_1
XFILLER_200_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21619_ _21635_/A vssd1 vssd1 vccd1 vccd1 _21619_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_540 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25387_ _27733_/Q input44/X _25391_/S vssd1 vssd1 vccd1 vccd1 _25388_/A sky130_fd_sc_hd__mux2_1
X_22599_ _22593_/X _22594_/X _22595_/X _22596_/X _22597_/X _22598_/X vssd1 vssd1 vccd1
+ vccd1 _22600_/A sky130_fd_sc_hd__mux4_1
XFILLER_127_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27126_ _27126_/CLK _27126_/D vssd1 vssd1 vccd1 vccd1 _27126_/Q sky130_fd_sc_hd__dfxtp_1
X_15140_ _26384_/Q _13350_/X _15140_/S vssd1 vssd1 vccd1 vccd1 _15141_/A sky130_fd_sc_hd__mux2_1
X_24338_ _24338_/A vssd1 vssd1 vccd1 vccd1 _27452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15071_ _14743_/X _26415_/Q _15079_/S vssd1 vssd1 vccd1 vccd1 _15072_/A sky130_fd_sc_hd__mux2_1
X_27057_ _23004_/X _27057_/D vssd1 vssd1 vccd1 vccd1 _27057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24269_ _24279_/A vssd1 vssd1 vccd1 vccd1 _24269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _26789_/Q _14005_/X _14019_/X _14021_/Y vssd1 vssd1 vccd1 vccd1 _26789_/D
+ sky130_fd_sc_hd__a31o_1
X_26008_ _27420_/CLK _26008_/D vssd1 vssd1 vccd1 vccd1 _26008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18830_ _18897_/A vssd1 vssd1 vccd1 vccd1 _19287_/A sky130_fd_sc_hd__buf_2
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18761_ _26041_/Q _17775_/X _18761_/S vssd1 vssd1 vccd1 vccd1 _18762_/A sky130_fd_sc_hd__mux2_1
X_15973_ _15973_/A vssd1 vssd1 vccd1 vccd1 _15973_/Y sky130_fd_sc_hd__inv_2
X_27959_ _27959_/A _15915_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17712_ _27419_/Q vssd1 vssd1 vccd1 vccd1 _17712_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14924_ _14924_/A vssd1 vssd1 vccd1 vccd1 _26473_/D sky130_fd_sc_hd__clkbuf_1
X_18692_ _18748_/A vssd1 vssd1 vccd1 vccd1 _18761_/S sky130_fd_sc_hd__buf_2
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17643_ _17482_/X _25893_/Q _17645_/S vssd1 vssd1 vccd1 vccd1 _17644_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14855_ _26503_/Q _13379_/X _14857_/S vssd1 vssd1 vccd1 vccd1 _14856_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13806_ _13844_/A vssd1 vssd1 vccd1 vccd1 _13806_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17574_ _17574_/A vssd1 vssd1 vccd1 vccd1 _25862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14786_ _14785_/X _26530_/Q _14789_/S vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16525_ _16824_/A _16257_/A _16292_/C _16292_/D _16106_/A vssd1 vssd1 vccd1 vccd1
+ _16526_/B sky130_fd_sc_hd__o41a_1
X_19313_ _19313_/A _19313_/B vssd1 vssd1 vccd1 vccd1 _19314_/A sky130_fd_sc_hd__and2_1
XFILLER_189_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13737_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19244_ _19241_/X _19243_/X _19334_/S vssd1 vssd1 vccd1 vccd1 _19244_/X sky130_fd_sc_hd__mux2_1
X_16456_ _16768_/B _16469_/B vssd1 vssd1 vccd1 vccd1 _16610_/A sky130_fd_sc_hd__xor2_1
X_13668_ _13938_/A _13670_/B vssd1 vssd1 vccd1 vccd1 _13668_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15407_ _15407_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15464_/A sky130_fd_sc_hd__nor2_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19175_ _19222_/A _19175_/B _19175_/C vssd1 vssd1 vccd1 vccd1 _19176_/A sky130_fd_sc_hd__and3_1
X_16387_ _16747_/B vssd1 vssd1 vccd1 vccd1 _16742_/A sky130_fd_sc_hd__clkbuf_2
X_13599_ _13639_/A vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18126_ _18425_/A vssd1 vssd1 vccd1 vccd1 _18126_/X sky130_fd_sc_hd__clkbuf_2
X_15338_ _14709_/X _26297_/Q _15346_/S vssd1 vssd1 vccd1 vccd1 _15339_/A sky130_fd_sc_hd__mux2_1
XFILLER_200_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18057_ _18479_/A vssd1 vssd1 vccd1 vccd1 _18057_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_0 _20349_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15269_ _26327_/Q _13328_/X _15273_/S vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ input8/X input7/X vssd1 vssd1 vccd1 vccd1 _23507_/A sky130_fd_sc_hd__nand2_4
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18959_ _18954_/X _18956_/X _18958_/X vssd1 vssd1 vccd1 vccd1 _18959_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21970_ _21986_/A vssd1 vssd1 vccd1 vccd1 _21970_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20921_ _20953_/A vssd1 vssd1 vccd1 vccd1 _20921_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23640_ _23638_/X _25733_/B _23640_/C vssd1 vssd1 vccd1 vccd1 _23641_/A sky130_fd_sc_hd__and3b_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20852_ _20852_/A vssd1 vssd1 vccd1 vccd1 _20852_/X sky130_fd_sc_hd__clkbuf_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23571_ _23577_/A _23571_/B vssd1 vssd1 vccd1 vccd1 _23572_/A sky130_fd_sc_hd__and2_1
XFILLER_23_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20783_ _20783_/A vssd1 vssd1 vccd1 vccd1 _20783_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25310_ _25310_/A _27512_/Q vssd1 vssd1 vccd1 vccd1 _25329_/C sky130_fd_sc_hd__xnor2_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22522_ _22522_/A vssd1 vssd1 vccd1 vccd1 _22522_/X sky130_fd_sc_hd__clkbuf_1
X_26290_ _20325_/X _26290_/D vssd1 vssd1 vccd1 vccd1 _26290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25241_ _25241_/A _25241_/B vssd1 vssd1 vccd1 vccd1 _25266_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22453_ _22453_/A vssd1 vssd1 vccd1 vccd1 _22520_/A sky130_fd_sc_hd__buf_2
XFILLER_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21404_ _21404_/A vssd1 vssd1 vccd1 vccd1 _21404_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25172_ _25164_/A _25171_/Y _25164_/B _25162_/A vssd1 vssd1 vccd1 vccd1 _25173_/B
+ sky130_fd_sc_hd__o31a_1
X_22384_ _22384_/A vssd1 vssd1 vccd1 vccd1 _22384_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24123_ _24123_/A vssd1 vssd1 vccd1 vccd1 _27335_/D sky130_fd_sc_hd__clkbuf_1
X_21335_ _21322_/X _21324_/X _21326_/X _21328_/X _21329_/X _21330_/X vssd1 vssd1 vccd1
+ vccd1 _21336_/A sky130_fd_sc_hd__mux4_1
XFILLER_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24054_ _24054_/A vssd1 vssd1 vccd1 vccd1 _27304_/D sky130_fd_sc_hd__clkbuf_1
X_21266_ _21266_/A vssd1 vssd1 vccd1 vccd1 _21266_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23005_ _22993_/X _22994_/X _22995_/X _22996_/X _22997_/X _22998_/X vssd1 vssd1 vccd1
+ vccd1 _23006_/A sky130_fd_sc_hd__mux4_1
X_20217_ _20249_/A vssd1 vssd1 vccd1 vccd1 _20217_/X sky130_fd_sc_hd__clkbuf_1
X_21197_ _21213_/A vssd1 vssd1 vccd1 vccd1 _21197_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27813_ _25698_/X _27813_/D vssd1 vssd1 vccd1 vccd1 _27813_/Q sky130_fd_sc_hd__dfxtp_1
X_20148_ _20164_/A vssd1 vssd1 vccd1 vccd1 _20148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12970_ _27812_/Q _12976_/B vssd1 vssd1 vccd1 vccd1 _12971_/A sky130_fd_sc_hd__and2_1
X_27744_ _27744_/CLK _27744_/D vssd1 vssd1 vccd1 vccd1 _27744_/Q sky130_fd_sc_hd__dfxtp_1
X_20079_ _20079_/A vssd1 vssd1 vccd1 vccd1 _20079_/X sky130_fd_sc_hd__clkbuf_1
X_24956_ _24960_/B _24956_/B vssd1 vssd1 vccd1 vccd1 _24957_/B sky130_fd_sc_hd__or2_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23907_ _24001_/A vssd1 vssd1 vccd1 vccd1 _23907_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27675_ _27675_/CLK _27675_/D vssd1 vssd1 vccd1 vccd1 _27966_/A sky130_fd_sc_hd__dfxtp_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24887_ _27767_/Q _24887_/B vssd1 vssd1 vccd1 vccd1 _24888_/B sky130_fd_sc_hd__nor2_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26626_ _21506_/X _26626_/D vssd1 vssd1 vccd1 vccd1 _26626_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14693_/A vssd1 vssd1 vccd1 vccd1 _14640_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23838_ _27074_/Q _27106_/Q _23845_/S vssd1 vssd1 vccd1 vccd1 _23838_/X sky130_fd_sc_hd__mux2_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _15732_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14571_/Y sky130_fd_sc_hd__nor2_1
X_26557_ _21264_/X _26557_/D vssd1 vssd1 vccd1 vccd1 _26557_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23769_ _23740_/X _23759_/X _23766_/X _23768_/X vssd1 vssd1 vccd1 vccd1 _27271_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16310_ _16310_/A vssd1 vssd1 vccd1 vccd1 _16412_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13522_ _13908_/A _13542_/B vssd1 vssd1 vccd1 vccd1 _13522_/Y sky130_fd_sc_hd__nor2_1
X_25508_ _24765_/A _25504_/X _25505_/Y _25507_/X _25497_/X vssd1 vssd1 vccd1 vccd1
+ _27765_/D sky130_fd_sc_hd__a221oi_1
XFILLER_201_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17290_ _17277_/X _17290_/B vssd1 vssd1 vccd1 vccd1 _17290_/X sky130_fd_sc_hd__and2b_1
XFILLER_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26488_ _21020_/X _26488_/D vssd1 vssd1 vccd1 vccd1 _26488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16241_ _27388_/Q _16132_/A _16137_/A _26054_/Q _16240_/X vssd1 vssd1 vccd1 vccd1
+ _24284_/A sky130_fd_sc_hd__a221o_1
X_13453_ _14433_/A vssd1 vssd1 vccd1 vccd1 _13870_/A sky130_fd_sc_hd__clkbuf_2
X_25439_ _25582_/A vssd1 vssd1 vccd1 vccd1 _25552_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_573 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16172_ _27576_/Q vssd1 vssd1 vccd1 vccd1 _16172_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_154_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ _13384_/A vssd1 vssd1 vccd1 vccd1 _26982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27109_ _27109_/CLK _27109_/D vssd1 vssd1 vccd1 vccd1 _27109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15123_ _26392_/Q _13325_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15124_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19931_ _19931_/A vssd1 vssd1 vccd1 vccd1 _19931_/X sky130_fd_sc_hd__clkbuf_1
X_15054_ _15054_/A vssd1 vssd1 vccd1 vccd1 _26423_/D sky130_fd_sc_hd__clkbuf_1
X_14005_ _14005_/A vssd1 vssd1 vccd1 vccd1 _14005_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19862_ _19850_/X _19851_/X _19852_/X _19853_/X _19854_/X _19855_/X vssd1 vssd1 vccd1
+ vccd1 _19863_/A sky130_fd_sc_hd__mux4_1
XFILLER_1_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18813_ _27600_/Q vssd1 vssd1 vccd1 vccd1 _18929_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19793_ _19793_/A vssd1 vssd1 vccd1 vccd1 _19793_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18744_ _26033_/Q _17750_/X _18746_/S vssd1 vssd1 vccd1 vccd1 _18745_/A sky130_fd_sc_hd__mux2_1
X_15956_ _15956_/A vssd1 vssd1 vccd1 vccd1 _15961_/A sky130_fd_sc_hd__buf_2
XFILLER_37_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14907_ _14740_/X _26480_/Q _14907_/S vssd1 vssd1 vccd1 vccd1 _14908_/A sky130_fd_sc_hd__mux2_1
X_18675_ _18675_/A vssd1 vssd1 vccd1 vccd1 _26002_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15887_ _15887_/A vssd1 vssd1 vccd1 vccd1 _15887_/Y sky130_fd_sc_hd__inv_2
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17626_ _17456_/X _25885_/Q _17634_/S vssd1 vssd1 vccd1 vccd1 _17627_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14838_ _26511_/Q _13353_/X _14846_/S vssd1 vssd1 vccd1 vccd1 _14839_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17557_ _17557_/A vssd1 vssd1 vccd1 vccd1 _25854_/D sky130_fd_sc_hd__clkbuf_1
X_14769_ _14769_/A vssd1 vssd1 vccd1 vccd1 _14769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _16508_/A _16508_/B vssd1 vssd1 vccd1 vccd1 _16508_/Y sky130_fd_sc_hd__nor2_1
X_17488_ _27428_/Q vssd1 vssd1 vccd1 vccd1 _17488_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19227_ _19227_/A vssd1 vssd1 vccd1 vccd1 _19227_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ _16772_/A _16256_/B _16767_/A _16486_/A vssd1 vssd1 vccd1 vccd1 _16440_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_158_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19158_ _19431_/A vssd1 vssd1 vccd1 vccd1 _19158_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_192_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18109_ _18057_/X _18105_/X _18108_/X _18062_/X vssd1 vssd1 vccd1 vccd1 _18109_/X
+ sky130_fd_sc_hd__o211a_1
X_19089_ _19387_/A vssd1 vssd1 vccd1 vccd1 _19089_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21120_ _21120_/A vssd1 vssd1 vccd1 vccd1 _21120_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21051_ _21039_/X _21040_/X _21041_/X _21042_/X _21044_/X _21046_/X vssd1 vssd1 vccd1
+ vccd1 _21052_/A sky130_fd_sc_hd__mux4_1
XFILLER_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20002_ _19988_/X _19989_/X _19990_/X _19991_/X _19994_/X _19997_/X vssd1 vssd1 vccd1
+ vccd1 _20003_/A sky130_fd_sc_hd__mux4_1
XFILLER_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24810_ _24960_/A vssd1 vssd1 vccd1 vccd1 _24811_/A sky130_fd_sc_hd__inv_2
X_25790_ _17501_/X _27850_/Q _25790_/S vssd1 vssd1 vccd1 vccd1 _25791_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24741_ _27612_/Q _24727_/X _24740_/Y _24729_/X vssd1 vssd1 vccd1 vccd1 _27612_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21953_ _21985_/A vssd1 vssd1 vccd1 vccd1 _21953_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20904_ _20904_/A vssd1 vssd1 vccd1 vccd1 _20904_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27460_ _27562_/CLK _27460_/D vssd1 vssd1 vccd1 vccd1 _27460_/Q sky130_fd_sc_hd__dfxtp_1
X_24672_ _27587_/Q _24660_/X _24671_/X _24663_/X vssd1 vssd1 vccd1 vccd1 _27587_/D
+ sky130_fd_sc_hd__o211a_1
X_21884_ _21900_/A vssd1 vssd1 vccd1 vccd1 _21884_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26411_ _20747_/X _26411_/D vssd1 vssd1 vccd1 vccd1 _26411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23623_ _27784_/Q _27226_/Q _23623_/S vssd1 vssd1 vccd1 vccd1 _23624_/B sky130_fd_sc_hd__mux2_1
X_20835_ _20867_/A vssd1 vssd1 vccd1 vccd1 _20835_/X sky130_fd_sc_hd__clkbuf_1
X_27391_ _27394_/CLK _27391_/D vssd1 vssd1 vccd1 vccd1 _27391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26342_ _20507_/X _26342_/D vssd1 vssd1 vccd1 vccd1 _26342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23554_ _23560_/A _23554_/B vssd1 vssd1 vccd1 vccd1 _23555_/A sky130_fd_sc_hd__and2_1
X_20766_ _20754_/X _20755_/X _20756_/X _20757_/X _20758_/X _20759_/X vssd1 vssd1 vccd1
+ vccd1 _20767_/A sky130_fd_sc_hd__mux4_1
XFILLER_74_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22505_ _22521_/A vssd1 vssd1 vccd1 vccd1 _22505_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_126_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26273_ _20263_/X _26273_/D vssd1 vssd1 vccd1 vccd1 _26273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_493 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23485_ _23485_/A vssd1 vssd1 vccd1 vccd1 _23495_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_168_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20697_ _20697_/A vssd1 vssd1 vccd1 vccd1 _20697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28012_ _28012_/A _15975_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_25224_ _25309_/A vssd1 vssd1 vccd1 vccd1 _25261_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_22436_ _22436_/A vssd1 vssd1 vccd1 vccd1 _22436_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1065 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25155_ _25155_/A _25164_/A vssd1 vssd1 vccd1 vccd1 _25157_/A sky130_fd_sc_hd__nor2_1
XFILLER_184_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22367_ _22453_/A vssd1 vssd1 vccd1 vccd1 _22434_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24106_ _27401_/Q _24106_/B vssd1 vssd1 vccd1 vccd1 _24107_/A sky130_fd_sc_hd__and2_1
X_21318_ _21318_/A vssd1 vssd1 vccd1 vccd1 _21318_/X sky130_fd_sc_hd__clkbuf_1
X_25086_ _25925_/Q _25991_/Q _25824_/Q _26023_/Q _25052_/X _25070_/X vssd1 vssd1 vccd1
+ vccd1 _25086_/X sky130_fd_sc_hd__mux4_1
X_22298_ _22298_/A vssd1 vssd1 vccd1 vccd1 _22298_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24037_ _25942_/Q _26008_/Q _25841_/Q _26040_/Q _23777_/A _23744_/A vssd1 vssd1 vccd1
+ vccd1 _24037_/X sky130_fd_sc_hd__mux4_1
X_21249_ _21231_/X _21234_/X _21237_/X _21240_/X _21241_/X _21242_/X vssd1 vssd1 vccd1
+ vccd1 _21250_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15810_ _13122_/X _26094_/Q _15816_/S vssd1 vssd1 vccd1 vccd1 _15811_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16790_ _16790_/A _16790_/B vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__xnor2_1
XFILLER_120_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25988_ _27140_/CLK _25988_/D vssd1 vssd1 vccd1 vccd1 _25988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ _15741_/A _15745_/B vssd1 vssd1 vccd1 vccd1 _15741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _12953_/A vssd1 vssd1 vccd1 vccd1 _27819_/D sky130_fd_sc_hd__clkbuf_1
X_27727_ _27729_/CLK _27727_/D vssd1 vssd1 vccd1 vccd1 _27727_/Q sky130_fd_sc_hd__dfxtp_1
X_24939_ _27664_/Q _24935_/X _24937_/Y _24938_/X vssd1 vssd1 vccd1 vccd1 _27664_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15672_ _13179_/X _26148_/Q _15678_/S vssd1 vssd1 vccd1 vccd1 _15673_/A sky130_fd_sc_hd__mux2_1
X_18460_ _18437_/X _18459_/X _18326_/X vssd1 vssd1 vccd1 vccd1 _18460_/X sky130_fd_sc_hd__o21a_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 _14788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27658_ _27658_/CLK _27658_/D vssd1 vssd1 vccd1 vccd1 _27658_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _25358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14707_/B sky130_fd_sc_hd__clkbuf_2
X_17411_ _27403_/Q _27402_/Q _27401_/Q _27400_/Q vssd1 vssd1 vccd1 vccd1 _17413_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA_242 _25639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26609_ _21442_/X _26609_/D vssd1 vssd1 vccd1 vccd1 _26609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_253 _27594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18391_ _18279_/X _18390_/X _18326_/X vssd1 vssd1 vccd1 vccd1 _18391_/X sky130_fd_sc_hd__o21a_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _25925_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27589_ _27589_/CLK _27589_/D vssd1 vssd1 vccd1 vccd1 _27589_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_286 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ input37/X vssd1 vssd1 vccd1 vccd1 _17342_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14554_ _15714_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14554_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_297 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13553_/A vssd1 vssd1 vccd1 vccd1 _13505_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17273_ _17271_/X _17272_/X _17296_/S vssd1 vssd1 vccd1 vccd1 _17273_/X sky130_fd_sc_hd__mux2_1
X_14485_ _16243_/A vssd1 vssd1 vccd1 vccd1 _15749_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_202_797 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16224_ _16224_/A _16224_/B _16235_/C vssd1 vssd1 vccd1 vccd1 _16224_/X sky130_fd_sc_hd__and3_1
X_19012_ _19012_/A vssd1 vssd1 vccd1 vccd1 _26048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13436_ _27365_/Q _13063_/X _13064_/X _27333_/Q _13056_/X vssd1 vssd1 vccd1 vccd1
+ _16099_/A sky130_fd_sc_hd__a221oi_4
XFILLER_174_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16155_ _16110_/A _24300_/A _16648_/A vssd1 vssd1 vccd1 vccd1 _16805_/A sky130_fd_sc_hd__o21ai_1
XFILLER_154_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13367_ _26987_/Q _13366_/X _13367_/S vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _14795_/X _26399_/Q _15112_/S vssd1 vssd1 vccd1 vccd1 _15107_/A sky130_fd_sc_hd__mux2_1
X_16086_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16650_/A sky130_fd_sc_hd__clkbuf_2
X_13298_ _27011_/Q _13184_/X _13302_/S vssd1 vssd1 vccd1 vccd1 _13299_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15037_ _26429_/Q _15028_/X _15029_/X _15036_/Y vssd1 vssd1 vccd1 vccd1 _26429_/D
+ sky130_fd_sc_hd__a31o_1
X_19914_ _19898_/X _19899_/X _19900_/X _19901_/X _19903_/X _19905_/X vssd1 vssd1 vccd1
+ vccd1 _19915_/A sky130_fd_sc_hd__mux4_1
X_19845_ _19845_/A vssd1 vssd1 vccd1 vccd1 _19845_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19776_ _19764_/X _19765_/X _19766_/X _19767_/X _19768_/X _19769_/X vssd1 vssd1 vccd1
+ vccd1 _19777_/A sky130_fd_sc_hd__mux4_1
XFILLER_84_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16988_ input36/X vssd1 vssd1 vccd1 vccd1 _17252_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18727_ _26025_/Q _17724_/X _18735_/S vssd1 vssd1 vccd1 vccd1 _18728_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15939_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18658_ _18658_/A vssd1 vssd1 vccd1 vccd1 _25994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17609_ _17609_/A vssd1 vssd1 vccd1 vccd1 _25877_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18589_ _24828_/A _25474_/A vssd1 vssd1 vccd1 vccd1 _18589_/X sky130_fd_sc_hd__or2_1
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20620_ _20706_/A vssd1 vssd1 vccd1 vccd1 _20686_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20551_ _20599_/A vssd1 vssd1 vccd1 vccd1 _20551_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23270_ _23254_/Y input69/X _23266_/Y input55/X _23269_/X vssd1 vssd1 vccd1 vccd1
+ _23275_/C sky130_fd_sc_hd__o221ai_1
XFILLER_158_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20482_ _20514_/A vssd1 vssd1 vccd1 vccd1 _20482_/X sky130_fd_sc_hd__clkbuf_1
X_22221_ _22213_/X _22214_/X _22215_/X _22216_/X _22217_/X _22218_/X vssd1 vssd1 vccd1
+ vccd1 _22222_/A sky130_fd_sc_hd__mux4_1
XFILLER_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22152_ _22152_/A vssd1 vssd1 vccd1 vccd1 _22152_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21103_ _21093_/X _21094_/X _21095_/X _21096_/X _21097_/X _21098_/X vssd1 vssd1 vccd1
+ vccd1 _21104_/A sky130_fd_sc_hd__mux4_1
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22083_ _22083_/A vssd1 vssd1 vccd1 vccd1 _22083_/X sky130_fd_sc_hd__clkbuf_1
X_26960_ _22672_/X _26960_/D vssd1 vssd1 vccd1 vccd1 _26960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21034_ _21034_/A vssd1 vssd1 vccd1 vccd1 _21034_/X sky130_fd_sc_hd__clkbuf_1
X_25911_ _27348_/CLK _25911_/D vssd1 vssd1 vccd1 vccd1 _25911_/Q sky130_fd_sc_hd__dfxtp_1
X_26891_ _22426_/X _26891_/D vssd1 vssd1 vccd1 vccd1 _26891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25842_ _27096_/CLK _25842_/D vssd1 vssd1 vccd1 vccd1 _25842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25773_ _17476_/X _27842_/Q _25779_/S vssd1 vssd1 vccd1 vccd1 _25774_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22985_ _22974_/X _22976_/X _22978_/X _22980_/X _22981_/X _22982_/X vssd1 vssd1 vccd1
+ vccd1 _22986_/A sky130_fd_sc_hd__mux4_1
XFILLER_16_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24724_ _27606_/Q _24714_/X _24723_/X _24717_/X vssd1 vssd1 vccd1 vccd1 _27606_/D
+ sky130_fd_sc_hd__o211a_1
X_27512_ _27515_/CLK _27512_/D vssd1 vssd1 vccd1 vccd1 _27512_/Q sky130_fd_sc_hd__dfxtp_1
X_21936_ _22000_/A vssd1 vssd1 vccd1 vccd1 _21936_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27443_ _27443_/CLK _27443_/D vssd1 vssd1 vccd1 vccd1 _27443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24655_ _27580_/Q _24643_/X _24654_/X _24650_/X vssd1 vssd1 vccd1 vccd1 _27580_/D
+ sky130_fd_sc_hd__o211a_1
X_21867_ _21899_/A vssd1 vssd1 vccd1 vccd1 _21867_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23606_ _23606_/A vssd1 vssd1 vccd1 vccd1 _27221_/D sky130_fd_sc_hd__clkbuf_1
X_20818_ _20866_/A vssd1 vssd1 vccd1 vccd1 _20818_/X sky130_fd_sc_hd__clkbuf_1
X_27374_ _27477_/CLK _27374_/D vssd1 vssd1 vccd1 vccd1 _27374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24586_ _24586_/A vssd1 vssd1 vccd1 vccd1 _27553_/D sky130_fd_sc_hd__clkbuf_1
X_21798_ _21814_/A vssd1 vssd1 vccd1 vccd1 _21798_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26325_ _20455_/X _26325_/D vssd1 vssd1 vccd1 vccd1 _26325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23537_ _23543_/A _23537_/B vssd1 vssd1 vccd1 vccd1 _23538_/A sky130_fd_sc_hd__and2_1
X_20749_ _20749_/A vssd1 vssd1 vccd1 vccd1 _20749_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_796 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14270_ _14296_/A vssd1 vssd1 vccd1 vccd1 _14270_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_26256_ _20209_/X _26256_/D vssd1 vssd1 vccd1 vccd1 _26256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23468_ input18/X _23455_/X _23467_/X _23461_/X vssd1 vssd1 vccd1 vccd1 _27180_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25207_ _27701_/Q _25184_/X _25206_/Y _25175_/X vssd1 vssd1 vccd1 vccd1 _27701_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_659 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13221_ _16197_/A vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__buf_2
XFILLER_100_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22419_ _22435_/A vssd1 vssd1 vccd1 vccd1 _22419_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26187_ _19967_/X _26187_/D vssd1 vssd1 vccd1 vccd1 _26187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23399_ _24752_/A _27240_/Q _27252_/Q _24782_/A _23398_/X vssd1 vssd1 vccd1 vccd1
+ _23409_/B sky130_fd_sc_hd__o221ai_1
XFILLER_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25138_ _25138_/A _25138_/B vssd1 vssd1 vccd1 vccd1 _25139_/B sky130_fd_sc_hd__xor2_1
X_13152_ _13152_/A vssd1 vssd1 vccd1 vccd1 _27049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_865 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25069_ _27837_/Q _27141_/Q _25886_/Q _25854_/Q _25061_/X _25035_/X vssd1 vssd1 vccd1
+ vccd1 _25069_/X sky130_fd_sc_hd__mux4_1
X_13083_ _27297_/Q _13109_/B vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__and2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17960_ _26142_/Q _26078_/Q _27006_/Q _26974_/Q _17870_/X _17959_/X vssd1 vssd1 vccd1
+ vccd1 _17961_/A sky130_fd_sc_hd__mux4_1
X_16911_ _16911_/A _16911_/B vssd1 vssd1 vccd1 vccd1 _16911_/Y sky130_fd_sc_hd__xnor2_1
X_17891_ _26812_/Q _26780_/Q _26748_/Q _26716_/Q _17863_/X _17890_/X vssd1 vssd1 vccd1
+ vccd1 _17891_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19630_ _19630_/A vssd1 vssd1 vccd1 vccd1 _19630_/X sky130_fd_sc_hd__clkbuf_1
X_16842_ _16864_/A _16842_/B vssd1 vssd1 vccd1 vccd1 _16843_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19561_ _26297_/Q _26265_/Q _26233_/Q _26201_/Q _18908_/X _19486_/X vssd1 vssd1 vccd1
+ vccd1 _19561_/X sky130_fd_sc_hd__mux4_1
X_13985_ _14359_/A _13992_/B vssd1 vssd1 vccd1 vccd1 _13985_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16773_ _16722_/X _16721_/A _16786_/A vssd1 vssd1 vccd1 vccd1 _16785_/A sky130_fd_sc_hd__a21oi_1
XFILLER_168_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18512_ _27821_/Q _26582_/Q _26454_/Q _26134_/Q _17899_/X _17901_/X vssd1 vssd1 vccd1
+ vccd1 _18512_/X sky130_fd_sc_hd__mux4_1
X_15724_ _26129_/Q _15721_/X _15713_/X _15723_/Y vssd1 vssd1 vccd1 vccd1 _26129_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12936_ input2/X _27858_/Q vssd1 vssd1 vccd1 vccd1 _13244_/B sky130_fd_sc_hd__nor2_4
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19492_ _19492_/A vssd1 vssd1 vccd1 vccd1 _19565_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18443_ _18443_/A vssd1 vssd1 vccd1 vccd1 _18443_/X sky130_fd_sc_hd__clkbuf_2
X_15655_ _15655_/A vssd1 vssd1 vccd1 vccd1 _26156_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _15767_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14606_/Y sky130_fd_sc_hd__nor2_1
X_15586_ _15608_/A vssd1 vssd1 vccd1 vccd1 _15595_/S sky130_fd_sc_hd__clkbuf_2
X_18374_ _18398_/A _18374_/B _18374_/C vssd1 vssd1 vccd1 vccd1 _18375_/A sky130_fd_sc_hd__and3_1
XFILLER_15_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14552_/A vssd1 vssd1 vccd1 vccd1 _14542_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17325_ _17325_/A vssd1 vssd1 vccd1 vccd1 _17325_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_18_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14468_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14483_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17256_ _25831_/Q _26030_/Q _17280_/S vssd1 vssd1 vccd1 vccd1 _17256_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16207_ _27526_/Q _16172_/X vssd1 vssd1 vccd1 vccd1 _16207_/X sky130_fd_sc_hd__or2b_1
X_13419_ _13419_/A vssd1 vssd1 vccd1 vccd1 _26971_/D sky130_fd_sc_hd__clkbuf_1
X_17187_ input38/X vssd1 vssd1 vccd1 vccd1 _17235_/S sky130_fd_sc_hd__clkbuf_2
X_14399_ _14399_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14399_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _16287_/A _16298_/C vssd1 vssd1 vccd1 vccd1 _16138_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16069_ _16457_/B vssd1 vssd1 vccd1 vccd1 _16402_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19828_ _19812_/X _19813_/X _19814_/X _19815_/X _19817_/X _19819_/X vssd1 vssd1 vccd1
+ vccd1 _19829_/A sky130_fd_sc_hd__mux4_1
XFILLER_151_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19759_ _19759_/A vssd1 vssd1 vccd1 vccd1 _19759_/X sky130_fd_sc_hd__clkbuf_1
X_22770_ _22786_/A vssd1 vssd1 vccd1 vccd1 _22770_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21721_ _21737_/A vssd1 vssd1 vccd1 vccd1 _21721_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_24440_ _24440_/A vssd1 vssd1 vccd1 vccd1 _27497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21652_ _21725_/A vssd1 vssd1 vccd1 vccd1 _21652_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20603_ _20672_/A vssd1 vssd1 vccd1 vccd1 _20603_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24371_ _24371_/A vssd1 vssd1 vccd1 vccd1 _27467_/D sky130_fd_sc_hd__clkbuf_1
X_21583_ _21583_/A vssd1 vssd1 vccd1 vccd1 _21649_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26110_ _19701_/X _26110_/D vssd1 vssd1 vccd1 vccd1 _26110_/Q sky130_fd_sc_hd__dfxtp_1
X_23322_ _23322_/A _23322_/B vssd1 vssd1 vccd1 vccd1 _23416_/A sky130_fd_sc_hd__nor2_1
X_27090_ _27123_/CLK _27090_/D vssd1 vssd1 vccd1 vccd1 _27090_/Q sky130_fd_sc_hd__dfxtp_1
X_20534_ _20706_/A vssd1 vssd1 vccd1 vccd1 _20600_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26041_ _27096_/CLK _26041_/D vssd1 vssd1 vccd1 vccd1 _26041_/Q sky130_fd_sc_hd__dfxtp_1
X_23253_ _23253_/A vssd1 vssd1 vccd1 vccd1 _27161_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_788 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20465_ _20513_/A vssd1 vssd1 vccd1 vccd1 _20465_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22204_ _22204_/A vssd1 vssd1 vccd1 vccd1 _22204_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23184_ _23252_/S vssd1 vssd1 vccd1 vccd1 _23193_/S sky130_fd_sc_hd__clkbuf_2
X_20396_ _20412_/A vssd1 vssd1 vccd1 vccd1 _20396_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22135_ _22125_/X _22126_/X _22127_/X _22128_/X _22129_/X _22130_/X vssd1 vssd1 vccd1
+ vccd1 _22136_/A sky130_fd_sc_hd__mux4_1
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27992_ _27992_/A _15890_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
XFILLER_160_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_813 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22066_ _22066_/A vssd1 vssd1 vccd1 vccd1 _22066_/X sky130_fd_sc_hd__clkbuf_1
X_26943_ _22606_/X _26943_/D vssd1 vssd1 vccd1 vccd1 _26943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21017_ _21007_/X _21008_/X _21009_/X _21010_/X _21011_/X _21012_/X vssd1 vssd1 vccd1
+ vccd1 _21018_/A sky130_fd_sc_hd__mux4_1
XFILLER_102_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26874_ _22364_/X _26874_/D vssd1 vssd1 vccd1 vccd1 _26874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25825_ _27081_/CLK _25825_/D vssd1 vssd1 vccd1 vccd1 _25825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ _13861_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13770_/Y sky130_fd_sc_hd__nor2_1
X_25756_ _25756_/A vssd1 vssd1 vccd1 vccd1 _27834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22968_ _22968_/A vssd1 vssd1 vccd1 vccd1 _22968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21919_ _21911_/X _21912_/X _21913_/X _21914_/X _21916_/X _21918_/X vssd1 vssd1 vccd1
+ vccd1 _21920_/A sky130_fd_sc_hd__mux4_1
X_24707_ _27184_/Q _24711_/B vssd1 vssd1 vccd1 vccd1 _24707_/X sky130_fd_sc_hd__or2_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25687_ _25673_/X _25674_/X _25675_/X _25676_/X _25677_/X _25678_/X vssd1 vssd1 vccd1
+ vccd1 _25688_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22899_ _22888_/X _22890_/X _22892_/X _22894_/X _22895_/X _22896_/X vssd1 vssd1 vccd1
+ vccd1 _22900_/A sky130_fd_sc_hd__mux4_1
X_15440_ _26251_/Q _13366_/X _15440_/S vssd1 vssd1 vccd1 vccd1 _15441_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27426_ _27427_/CLK _27426_/D vssd1 vssd1 vccd1 vccd1 _27426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24638_ _24638_/A _24638_/B vssd1 vssd1 vccd1 vccd1 _24639_/A sky130_fd_sc_hd__and2_1
XFILLER_130_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15371_ _14759_/X _26282_/Q _15379_/S vssd1 vssd1 vccd1 vccd1 _15372_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24569_ _24569_/A vssd1 vssd1 vccd1 vccd1 _27545_/D sky130_fd_sc_hd__clkbuf_1
X_27357_ _27357_/CLK _27357_/D vssd1 vssd1 vccd1 vccd1 _27357_/Q sky130_fd_sc_hd__dfxtp_2
X_14322_ _14365_/A vssd1 vssd1 vccd1 vccd1 _14322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17110_ _17057_/X _17109_/X _17098_/X vssd1 vssd1 vccd1 vccd1 _17110_/X sky130_fd_sc_hd__a21bo_1
XFILLER_196_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18090_ _26403_/Q _26371_/Q _26339_/Q _26307_/Q _17903_/X _17904_/X vssd1 vssd1 vccd1
+ vccd1 _18090_/X sky130_fd_sc_hd__mux4_1
X_26308_ _20389_/X _26308_/D vssd1 vssd1 vccd1 vccd1 _26308_/Q sky130_fd_sc_hd__dfxtp_1
X_27288_ _27288_/CLK _27288_/D vssd1 vssd1 vccd1 vccd1 _27288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17041_ _25915_/Q _25981_/Q _17071_/S vssd1 vssd1 vccd1 vccd1 _17042_/B sky130_fd_sc_hd__mux2_1
X_14253_ _26710_/Q _14238_/X _14242_/X _14252_/Y vssd1 vssd1 vccd1 vccd1 _26710_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26239_ _20145_/X _26239_/D vssd1 vssd1 vccd1 vccd1 _26239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13204_ _14791_/A vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14184_ _14361_/A _14187_/B vssd1 vssd1 vccd1 vccd1 _14184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13135_ _13135_/A vssd1 vssd1 vccd1 vccd1 _27052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _19473_/A vssd1 vssd1 vccd1 vccd1 _19107_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_673 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _27364_/Q _13063_/X _13064_/X _27332_/Q _13065_/X vssd1 vssd1 vccd1 vccd1
+ _14718_/A sky130_fd_sc_hd__a221o_2
X_17943_ _18418_/A vssd1 vssd1 vccd1 vccd1 _17943_/X sky130_fd_sc_hd__clkbuf_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater207 _25987_/CLK vssd1 vssd1 vccd1 vccd1 _25986_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater218 _27397_/CLK vssd1 vssd1 vccd1 vccd1 _27302_/CLK sky130_fd_sc_hd__clkbuf_1
X_17874_ _26267_/Q _26235_/Q _26203_/Q _26171_/Q _17873_/X _17835_/X vssd1 vssd1 vccd1
+ vccd1 _17874_/X sky130_fd_sc_hd__mux4_1
Xrepeater229 _26073_/CLK vssd1 vssd1 vccd1 vccd1 _26067_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19613_ _19605_/X _19606_/X _19607_/X _19608_/X _19609_/X _19610_/X vssd1 vssd1 vccd1
+ vccd1 _19614_/A sky130_fd_sc_hd__mux4_1
X_16825_ _16805_/Y _16823_/X _16824_/Y vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19544_ _19485_/X _19543_/X _19488_/X vssd1 vssd1 vccd1 vccd1 _19544_/X sky130_fd_sc_hd__o21a_1
X_16756_ _16756_/A _16756_/B vssd1 vssd1 vccd1 vccd1 _16756_/X sky130_fd_sc_hd__or2_1
XFILLER_81_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13968_ _26804_/Q _13949_/X _13965_/X _13967_/Y vssd1 vssd1 vccd1 vccd1 _26804_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ _15761_/A vssd1 vssd1 vccd1 vccd1 _15718_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19475_ _19534_/A _19475_/B vssd1 vssd1 vccd1 vccd1 _19475_/X sky130_fd_sc_hd__or2_1
X_12919_ input53/X input54/X input55/X input56/X vssd1 vssd1 vccd1 vccd1 _12921_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_62_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13899_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13899_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16687_ _16686_/A _16686_/B _16619_/A vssd1 vssd1 vccd1 vccd1 _16687_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18426_ _27817_/Q _26578_/Q _26450_/Q _26130_/Q _18401_/X _18425_/X vssd1 vssd1 vccd1
+ vccd1 _18426_/X sky130_fd_sc_hd__mux4_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15638_ _15638_/A vssd1 vssd1 vccd1 vccd1 _26164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18357_ _18355_/X _18356_/X _18378_/S vssd1 vssd1 vccd1 vccd1 _18357_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15569_ _26194_/Q _14734_/A _15573_/S vssd1 vssd1 vccd1 vccd1 _15570_/A sky130_fd_sc_hd__mux2_1
X_17308_ _27090_/Q _27122_/Q _17355_/S vssd1 vssd1 vccd1 vccd1 _17308_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18288_ _18288_/A vssd1 vssd1 vccd1 vccd1 _25961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17239_ _27845_/Q _27149_/Q _25894_/Q _25862_/Q _17203_/X _17191_/X vssd1 vssd1 vccd1
+ vccd1 _17239_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20250_ _20250_/A vssd1 vssd1 vccd1 vccd1 _20250_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20181_ _20248_/A vssd1 vssd1 vccd1 vccd1 _20181_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23940_ _23938_/X _23939_/X _23940_/S vssd1 vssd1 vccd1 vccd1 _23940_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23871_ _27077_/Q _23860_/X _23861_/X _27109_/Q _23862_/X vssd1 vssd1 vccd1 vccd1
+ _23871_/X sky130_fd_sc_hd__a221o_1
X_25610_ _24815_/A _18606_/X _25608_/X _25609_/Y _25592_/X vssd1 vssd1 vccd1 vccd1
+ _27783_/D sky130_fd_sc_hd__a221oi_1
XFILLER_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22822_ _22870_/A vssd1 vssd1 vccd1 vccd1 _22822_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26590_ _21380_/X _26590_/D vssd1 vssd1 vccd1 vccd1 _26590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25541_ _27707_/Q _25539_/X _25540_/X vssd1 vssd1 vccd1 vccd1 _25541_/Y sky130_fd_sc_hd__a21oi_1
X_22753_ _22785_/A vssd1 vssd1 vccd1 vccd1 _22753_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_825 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21704_ _21704_/A vssd1 vssd1 vccd1 vccd1 _21704_/X sky130_fd_sc_hd__clkbuf_1
X_25472_ _25470_/X _25158_/B _25471_/X _25452_/X vssd1 vssd1 vccd1 vccd1 _25472_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_198_869 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22684_ _22700_/A vssd1 vssd1 vccd1 vccd1 _22684_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27211_ _27211_/CLK _27211_/D vssd1 vssd1 vccd1 vccd1 _27211_/Q sky130_fd_sc_hd__dfxtp_1
X_24423_ _24423_/A vssd1 vssd1 vccd1 vccd1 _27490_/D sky130_fd_sc_hd__clkbuf_1
X_21635_ _21635_/A vssd1 vssd1 vccd1 vccd1 _21635_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27142_ _27142_/CLK _27142_/D vssd1 vssd1 vccd1 vccd1 _27142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24354_ _24354_/A vssd1 vssd1 vccd1 vccd1 _27459_/D sky130_fd_sc_hd__clkbuf_1
X_21566_ _21635_/A vssd1 vssd1 vccd1 vccd1 _21566_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23305_ input72/X vssd1 vssd1 vccd1 vccd1 _23305_/Y sky130_fd_sc_hd__inv_2
X_20517_ _20586_/A vssd1 vssd1 vccd1 vccd1 _20517_/X sky130_fd_sc_hd__clkbuf_2
X_27073_ _27103_/CLK _27073_/D vssd1 vssd1 vccd1 vccd1 _27073_/Q sky130_fd_sc_hd__dfxtp_1
X_24285_ _24285_/A vssd1 vssd1 vccd1 vccd1 _27420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21497_ _21583_/A vssd1 vssd1 vccd1 vccd1 _21563_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_153_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26024_ _26024_/CLK _26024_/D vssd1 vssd1 vccd1 vccd1 _26024_/Q sky130_fd_sc_hd__dfxtp_1
X_23236_ _23236_/A vssd1 vssd1 vccd1 vccd1 _27153_/D sky130_fd_sc_hd__clkbuf_1
X_20448_ _20706_/A vssd1 vssd1 vccd1 vccd1 _20514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23167_ _23167_/A vssd1 vssd1 vccd1 vccd1 _23176_/S sky130_fd_sc_hd__buf_2
X_20379_ _20427_/A vssd1 vssd1 vccd1 vccd1 _20379_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22118_ _22118_/A vssd1 vssd1 vccd1 vccd1 _22118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23098_ _23098_/A vssd1 vssd1 vccd1 vccd1 _27092_/D sky130_fd_sc_hd__clkbuf_1
X_27975_ _27975_/A _15910_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22049_ _22035_/X _22036_/X _22037_/X _22038_/X _22039_/X _22040_/X vssd1 vssd1 vccd1
+ vccd1 _22050_/A sky130_fd_sc_hd__mux4_1
X_26926_ _22554_/X _26926_/D vssd1 vssd1 vccd1 vccd1 _26926_/Q sky130_fd_sc_hd__dfxtp_1
X_14940_ _14788_/X _26465_/Q _14940_/S vssd1 vssd1 vccd1 vccd1 _14941_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_571 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26857_ _22310_/X _26857_/D vssd1 vssd1 vccd1 vccd1 _26857_/Q sky130_fd_sc_hd__dfxtp_1
X_14871_ _26496_/Q _13401_/X _14879_/S vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16610_ _16610_/A _16610_/B vssd1 vssd1 vccd1 vccd1 _16610_/X sky130_fd_sc_hd__xor2_1
X_13822_ _26853_/Q _13819_/X _13820_/X _13821_/Y vssd1 vssd1 vccd1 vccd1 _26853_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25808_ _25808_/A vssd1 vssd1 vccd1 vccd1 _25808_/X sky130_fd_sc_hd__clkbuf_1
X_17590_ _17590_/A vssd1 vssd1 vccd1 vccd1 _25869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26788_ _22064_/X _26788_/D vssd1 vssd1 vccd1 vccd1 _26788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13753_ _13934_/A _13759_/B vssd1 vssd1 vccd1 vccd1 _13753_/Y sky130_fd_sc_hd__nor2_1
X_16541_ _16616_/A _16616_/B vssd1 vssd1 vccd1 vccd1 _16885_/A sky130_fd_sc_hd__xor2_1
XFILLER_28_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25739_ _25739_/A vssd1 vssd1 vccd1 vccd1 _27826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19260_ _26155_/Q _26091_/Q _27019_/Q _26987_/Q _19165_/X _19188_/X vssd1 vssd1 vccd1
+ vccd1 _19261_/B sky130_fd_sc_hd__mux4_1
XFILLER_188_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13684_ _26903_/Q _13682_/X _13676_/X _13683_/Y vssd1 vssd1 vccd1 vccd1 _26903_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16472_ _16611_/B _16469_/B _16609_/A vssd1 vssd1 vccd1 vccd1 _16472_/X sky130_fd_sc_hd__o21ba_1
X_27961__447 vssd1 vssd1 vccd1 vccd1 _27961__447/HI _27961_/A sky130_fd_sc_hd__conb_1
X_18211_ _18483_/A vssd1 vssd1 vccd1 vccd1 _18211_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15423_ _26259_/Q _13341_/X _15429_/S vssd1 vssd1 vccd1 vccd1 _15424_/A sky130_fd_sc_hd__mux2_1
X_27409_ _27411_/CLK _27409_/D vssd1 vssd1 vccd1 vccd1 _27409_/Q sky130_fd_sc_hd__dfxtp_1
X_19191_ _19485_/A vssd1 vssd1 vccd1 vccd1 _19191_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18142_ _26533_/Q _26501_/Q _26469_/Q _27045_/Q _18117_/X _18141_/X vssd1 vssd1 vccd1
+ vccd1 _18142_/X sky130_fd_sc_hd__mux4_1
X_15354_ _15354_/A vssd1 vssd1 vccd1 vccd1 _26290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14305_ _14394_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14305_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18073_ _18418_/A vssd1 vssd1 vccd1 vccd1 _18073_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15285_ _15285_/A vssd1 vssd1 vccd1 vccd1 _26320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14236_ _15773_/A vssd1 vssd1 vccd1 vccd1 _14548_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17024_ _27067_/Q _27099_/Q _17047_/S vssd1 vssd1 vccd1 vccd1 _17024_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _14220_/A vssd1 vssd1 vccd1 vccd1 _14167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _27055_/Q _13116_/X _13140_/S vssd1 vssd1 vccd1 vccd1 _13119_/A sky130_fd_sc_hd__mux2_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14363_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14098_/Y sky130_fd_sc_hd__nor2_1
X_18975_ _27798_/Q _26559_/Q _26431_/Q _26111_/Q _18974_/X _18851_/X vssd1 vssd1 vccd1
+ vccd1 _18975_/X sky130_fd_sc_hd__mux4_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17926_ _17921_/X _17923_/X _18056_/S vssd1 vssd1 vccd1 vccd1 _17926_/X sky130_fd_sc_hd__mux2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _14885_/A _15695_/D vssd1 vssd1 vccd1 vccd1 _13205_/A sky130_fd_sc_hd__nor2_2
XFILLER_61_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17857_ _17828_/X _17839_/X _17852_/X _17854_/X _17856_/X vssd1 vssd1 vccd1 vccd1
+ _17858_/C sky130_fd_sc_hd__a221o_1
XFILLER_61_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16808_ _16808_/A _16808_/B vssd1 vssd1 vccd1 vccd1 _16811_/C sky130_fd_sc_hd__or2_1
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17788_ _17898_/A vssd1 vssd1 vccd1 vccd1 _18401_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19527_ _26423_/Q _26391_/Q _26359_/Q _26327_/Q _19465_/X _18795_/X vssd1 vssd1 vccd1
+ vccd1 _19527_/X sky130_fd_sc_hd__mux4_1
X_16739_ _16625_/A _16747_/A _16742_/A _16625_/B vssd1 vssd1 vccd1 vccd1 _16739_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_34_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19458_ _19456_/X _19457_/X _19480_/S vssd1 vssd1 vccd1 vccd1 _19458_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18409_ _26705_/Q _26673_/Q _26641_/Q _26609_/Q _18360_/X _18408_/X vssd1 vssd1 vccd1
+ vccd1 _18410_/A sky130_fd_sc_hd__mux4_2
XFILLER_14_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _26961_/Q _26929_/Q _26897_/Q _26865_/Q _19343_/X _19253_/X vssd1 vssd1 vccd1
+ vccd1 _19389_/X sky130_fd_sc_hd__mux4_1
XFILLER_194_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21420_ _21420_/A vssd1 vssd1 vccd1 vccd1 _21420_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21351_ _21341_/X _21342_/X _21343_/X _21344_/X _21345_/X _21346_/X vssd1 vssd1 vccd1
+ vccd1 _21352_/A sky130_fd_sc_hd__mux4_1
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20302_ _20334_/A vssd1 vssd1 vccd1 vccd1 _20302_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24070_ _27385_/Q _24072_/B vssd1 vssd1 vccd1 vccd1 _24071_/A sky130_fd_sc_hd__and2_1
X_21282_ _21282_/A vssd1 vssd1 vccd1 vccd1 _21282_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23021_ _23009_/X _23010_/X _23011_/X _23012_/X _23013_/X _23014_/X vssd1 vssd1 vccd1
+ vccd1 _23022_/A sky130_fd_sc_hd__mux4_1
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20233_ _20249_/A vssd1 vssd1 vccd1 vccd1 _20233_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20164_ _20164_/A vssd1 vssd1 vccd1 vccd1 _20164_/X sky130_fd_sc_hd__clkbuf_1
X_27760_ _27760_/CLK _27760_/D vssd1 vssd1 vccd1 vccd1 _27760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24972_ _25018_/A vssd1 vssd1 vccd1 vccd1 _24972_/X sky130_fd_sc_hd__buf_2
X_20095_ _20162_/A vssd1 vssd1 vccd1 vccd1 _20095_/X sky130_fd_sc_hd__clkbuf_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26711_ _21802_/X _26711_/D vssd1 vssd1 vccd1 vccd1 _26711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23923_ _23921_/X _23922_/X _23938_/S vssd1 vssd1 vccd1 vccd1 _23923_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27691_ _27693_/CLK _27691_/D vssd1 vssd1 vccd1 vccd1 _27691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26642_ _21556_/X _26642_/D vssd1 vssd1 vccd1 vccd1 _26642_/Q sky130_fd_sc_hd__dfxtp_1
X_23854_ _24045_/S vssd1 vssd1 vccd1 vccd1 _23891_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22805_ _22891_/A vssd1 vssd1 vccd1 vccd1 _22871_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26573_ _21318_/X _26573_/D vssd1 vssd1 vccd1 vccd1 _26573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23785_ _27829_/Q _27133_/Q _25878_/Q _25846_/Q _23777_/X _23744_/X vssd1 vssd1 vccd1
+ vccd1 _23785_/X sky130_fd_sc_hd__mux4_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20997_ _20991_/X _20992_/X _20993_/X _20994_/X _20995_/X _20996_/X vssd1 vssd1 vccd1
+ vccd1 _20998_/A sky130_fd_sc_hd__mux4_1
XFILLER_198_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25524_ _25524_/A vssd1 vssd1 vccd1 vccd1 _25524_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_22736_ _22784_/A vssd1 vssd1 vccd1 vccd1 _22736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25455_ _27693_/Q _25448_/X _25449_/X vssd1 vssd1 vccd1 vccd1 _25455_/Y sky130_fd_sc_hd__a21oi_1
X_22667_ _22699_/A vssd1 vssd1 vccd1 vccd1 _22667_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24406_ _24406_/A vssd1 vssd1 vccd1 vccd1 _27482_/D sky130_fd_sc_hd__clkbuf_1
X_21618_ _21650_/A vssd1 vssd1 vccd1 vccd1 _21618_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25386_ _25386_/A vssd1 vssd1 vccd1 vccd1 _27732_/D sky130_fd_sc_hd__clkbuf_1
X_22598_ _22598_/A vssd1 vssd1 vccd1 vccd1 _22598_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_27125_ _27125_/CLK _27125_/D vssd1 vssd1 vccd1 vccd1 _27125_/Q sky130_fd_sc_hd__dfxtp_1
X_24337_ _27552_/Q _24339_/B vssd1 vssd1 vccd1 vccd1 _24338_/A sky130_fd_sc_hd__and2_1
X_21549_ _21549_/A vssd1 vssd1 vccd1 vccd1 _21549_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15070_ _15116_/S vssd1 vssd1 vccd1 vccd1 _15079_/S sky130_fd_sc_hd__clkbuf_2
X_27056_ _23002_/X _27056_/D vssd1 vssd1 vccd1 vccd1 _27056_/Q sky130_fd_sc_hd__dfxtp_1
X_24268_ _24268_/A vssd1 vssd1 vccd1 vccd1 _27407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _14386_/A _14029_/B vssd1 vssd1 vccd1 vccd1 _14021_/Y sky130_fd_sc_hd__nor2_1
X_26007_ _26007_/CLK _26007_/D vssd1 vssd1 vccd1 vccd1 _26007_/Q sky130_fd_sc_hd__dfxtp_1
X_23219_ _23219_/A vssd1 vssd1 vccd1 vccd1 _27145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24199_ _24363_/A vssd1 vssd1 vccd1 vccd1 _24279_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18760_ _18760_/A vssd1 vssd1 vccd1 vccd1 _26040_/D sky130_fd_sc_hd__clkbuf_1
X_27958_ _27958_/A _15914_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
X_15972_ _15973_/A vssd1 vssd1 vccd1 vccd1 _15972_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17711_ _17711_/A vssd1 vssd1 vccd1 vccd1 _25922_/D sky130_fd_sc_hd__clkbuf_1
X_26909_ _22486_/X _26909_/D vssd1 vssd1 vccd1 vccd1 _26909_/Q sky130_fd_sc_hd__dfxtp_1
X_14923_ _14763_/X _26473_/Q _14929_/S vssd1 vssd1 vccd1 vccd1 _14924_/A sky130_fd_sc_hd__mux2_1
X_18691_ _18691_/A _18691_/B vssd1 vssd1 vccd1 vccd1 _18748_/A sky130_fd_sc_hd__nor2_2
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17642_ _17642_/A vssd1 vssd1 vccd1 vccd1 _25892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14854_ _14854_/A vssd1 vssd1 vccd1 vccd1 _26504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13805_ _26859_/Q _13793_/X _13794_/X _13804_/Y vssd1 vssd1 vccd1 vccd1 _26859_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_189_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17573_ _17485_/X _25862_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14785_ _14785_/A vssd1 vssd1 vccd1 vccd1 _14785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19312_ _19302_/X _19310_/X _19312_/S vssd1 vssd1 vccd1 vccd1 _19313_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16524_ _16036_/X _24301_/A _16648_/A vssd1 vssd1 vccd1 vccd1 _16908_/B sky130_fd_sc_hd__o21ai_4
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13736_ _26884_/Q _13724_/X _13732_/X _13735_/Y vssd1 vssd1 vccd1 vccd1 _26884_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19243_ _26538_/Q _26506_/Q _26474_/Q _27050_/Q _19242_/X _19148_/X vssd1 vssd1 vccd1
+ vccd1 _19243_/X sky130_fd_sc_hd__mux4_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16455_ _16783_/A _16455_/B vssd1 vssd1 vccd1 vccd1 _16469_/B sky130_fd_sc_hd__xnor2_2
XFILLER_143_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13667_ _26908_/Q _13665_/X _13656_/X _13666_/Y vssd1 vssd1 vccd1 vccd1 _26908_/D
+ sky130_fd_sc_hd__a31o_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15406_/A vssd1 vssd1 vccd1 vccd1 _26266_/D sky130_fd_sc_hd__clkbuf_1
X_19174_ _19167_/X _19169_/X _19173_/X _19151_/X _19105_/X vssd1 vssd1 vccd1 vccd1
+ _19175_/C sky130_fd_sc_hd__a221o_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _26934_/Q _13580_/X _13587_/X _13597_/Y vssd1 vssd1 vccd1 vccd1 _26934_/D
+ sky130_fd_sc_hd__a31o_1
X_16386_ _14791_/A _16384_/X _16375_/B _25950_/Q _16385_/Y vssd1 vssd1 vccd1 vccd1
+ _16747_/B sky130_fd_sc_hd__a221o_1
XFILLER_118_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18125_ _18125_/A vssd1 vssd1 vccd1 vccd1 _25954_/D sky130_fd_sc_hd__clkbuf_1
X_15337_ _15405_/S vssd1 vssd1 vccd1 vccd1 _15346_/S sky130_fd_sc_hd__buf_2
XFILLER_184_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18056_ _18054_/X _18055_/X _18056_/S vssd1 vssd1 vccd1 vccd1 _18056_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _20457_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _15268_/A vssd1 vssd1 vccd1 vccd1 _26328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17007_ _17003_/X _17005_/X _17048_/S vssd1 vssd1 vccd1 vccd1 _17007_/X sky130_fd_sc_hd__mux2_1
X_14219_ _26721_/Q _14212_/X _14207_/X _14218_/Y vssd1 vssd1 vccd1 vccd1 _26721_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15199_ _14721_/X _26358_/Q _15201_/S vssd1 vssd1 vccd1 vccd1 _15200_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18958_ _19488_/A vssd1 vssd1 vccd1 vccd1 _18958_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17909_ _26140_/Q _26076_/Q _27004_/Q _26972_/Q _17821_/X _24386_/A vssd1 vssd1 vccd1
+ vccd1 _17911_/A sky130_fd_sc_hd__mux4_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18889_ _26524_/Q _26492_/Q _26460_/Q _27036_/Q _18829_/X _18863_/X vssd1 vssd1 vccd1
+ vccd1 _18889_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20920_ _20920_/A vssd1 vssd1 vccd1 vccd1 _20920_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20851_ _20867_/A vssd1 vssd1 vccd1 vccd1 _20851_/X sky130_fd_sc_hd__clkbuf_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23570_ _27770_/Q _27212_/Q _23576_/S vssd1 vssd1 vccd1 vccd1 _23571_/B sky130_fd_sc_hd__mux2_1
XFILLER_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20782_ _20770_/X _20771_/X _20772_/X _20773_/X _20775_/X _20777_/X vssd1 vssd1 vccd1
+ vccd1 _20783_/A sky130_fd_sc_hd__mux4_1
XFILLER_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22521_ _22521_/A vssd1 vssd1 vccd1 vccd1 _22521_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25240_ _27536_/Q _27504_/Q vssd1 vssd1 vccd1 vccd1 _25241_/B sky130_fd_sc_hd__or2_1
X_22452_ _22519_/A vssd1 vssd1 vccd1 vccd1 _22452_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21403_ _21389_/X _21390_/X _21391_/X _21392_/X _21394_/X _21396_/X vssd1 vssd1 vccd1
+ vccd1 _21404_/A sky130_fd_sc_hd__mux4_1
X_25171_ _27526_/Q _27494_/Q vssd1 vssd1 vccd1 vccd1 _25171_/Y sky130_fd_sc_hd__nor2_1
X_22383_ _22366_/X _22368_/X _22370_/X _22372_/X _22373_/X _22374_/X vssd1 vssd1 vccd1
+ vccd1 _22384_/A sky130_fd_sc_hd__mux4_1
XFILLER_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24122_ _27440_/Q _24128_/B vssd1 vssd1 vccd1 vccd1 _24123_/A sky130_fd_sc_hd__and2_1
XFILLER_198_1173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21334_ _21334_/A vssd1 vssd1 vccd1 vccd1 _21334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24053_ _27377_/Q _24061_/B vssd1 vssd1 vccd1 vccd1 _24054_/A sky130_fd_sc_hd__and2_1
X_21265_ _21253_/X _21254_/X _21255_/X _21256_/X _21257_/X _21258_/X vssd1 vssd1 vccd1
+ vccd1 _21266_/A sky130_fd_sc_hd__mux4_1
XFILLER_117_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23004_ _23004_/A vssd1 vssd1 vccd1 vccd1 _23004_/X sky130_fd_sc_hd__clkbuf_1
X_20216_ _20248_/A vssd1 vssd1 vccd1 vccd1 _20216_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21196_ _21212_/A vssd1 vssd1 vccd1 vccd1 _21196_/X sky130_fd_sc_hd__clkbuf_1
X_27812_ _25696_/X _27812_/D vssd1 vssd1 vccd1 vccd1 _27812_/Q sky130_fd_sc_hd__dfxtp_1
X_20147_ _20163_/A vssd1 vssd1 vccd1 vccd1 _20147_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27743_ _27745_/CLK _27743_/D vssd1 vssd1 vccd1 vccd1 _27743_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _20078_/A vssd1 vssd1 vccd1 vccd1 _20078_/X sky130_fd_sc_hd__clkbuf_1
X_24955_ _24954_/B _24954_/C _25601_/A vssd1 vssd1 vccd1 vccd1 _24956_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23906_ _23902_/X _23904_/X _23940_/S vssd1 vssd1 vccd1 vccd1 _23906_/X sky130_fd_sc_hd__mux2_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27674_ _27674_/CLK _27674_/D vssd1 vssd1 vccd1 vccd1 _27965_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24886_ _27767_/Q _24887_/B vssd1 vssd1 vccd1 vccd1 _24896_/C sky130_fd_sc_hd__and2_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater390 _27222_/CLK vssd1 vssd1 vccd1 vccd1 _27196_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26625_ _21504_/X _26625_/D vssd1 vssd1 vccd1 vccd1 _26625_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23837_ _23834_/X _23836_/X _23844_/S vssd1 vssd1 vccd1 vccd1 _23837_/X sky130_fd_sc_hd__mux2_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _26606_/Q _14563_/X _14566_/X _14569_/Y vssd1 vssd1 vccd1 vccd1 _26606_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26556_ _21262_/X _26556_/D vssd1 vssd1 vccd1 vccd1 _26556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23768_ _23864_/A vssd1 vssd1 vccd1 vccd1 _23768_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_199_964 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13521_ _13546_/A vssd1 vssd1 vccd1 vccd1 _13542_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_25507_ _25500_/X _25206_/B _25506_/X _25483_/X vssd1 vssd1 vccd1 vccd1 _25507_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22719_ _22891_/A vssd1 vssd1 vccd1 vccd1 _22785_/A sky130_fd_sc_hd__buf_2
XFILLER_186_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23699_ _24925_/B _27254_/Q _23705_/S vssd1 vssd1 vccd1 vccd1 _23700_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26487_ _21018_/X _26487_/D vssd1 vssd1 vccd1 vccd1 _26487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_968 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _27362_/Q _13450_/X _13451_/X _27330_/Q _13075_/X vssd1 vssd1 vccd1 vccd1
+ _14433_/A sky130_fd_sc_hd__a221oi_4
X_16240_ _16240_/A _16249_/B _16240_/C vssd1 vssd1 vccd1 vccd1 _16240_/X sky130_fd_sc_hd__and3_1
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25438_ _25560_/A vssd1 vssd1 vccd1 vccd1 _25438_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25369_ _27725_/Q input67/X _25369_/S vssd1 vssd1 vccd1 vccd1 _25370_/A sky130_fd_sc_hd__mux2_1
X_13383_ _26982_/Q _13382_/X _13383_/S vssd1 vssd1 vccd1 vccd1 _13384_/A sky130_fd_sc_hd__mux2_1
X_16171_ _16034_/A _16166_/X _16168_/Y _16169_/X _16170_/X vssd1 vssd1 vccd1 vccd1
+ _16428_/A sky130_fd_sc_hd__o41a_1
XFILLER_182_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27108_ _27110_/CLK _27108_/D vssd1 vssd1 vccd1 vccd1 _27108_/Q sky130_fd_sc_hd__dfxtp_1
X_15122_ _15122_/A vssd1 vssd1 vccd1 vccd1 _26393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19930_ _19918_/X _19921_/X _19924_/X _19927_/X _19928_/X _19929_/X vssd1 vssd1 vccd1
+ vccd1 _19931_/A sky130_fd_sc_hd__mux4_1
X_15053_ _14718_/X _26423_/Q _15057_/S vssd1 vssd1 vccd1 vccd1 _15054_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27039_ _22938_/X _27039_/D vssd1 vssd1 vccd1 vccd1 _27039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14004_ _26794_/Q _13987_/X _14001_/X _14003_/Y vssd1 vssd1 vccd1 vccd1 _26794_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19861_ _19861_/A vssd1 vssd1 vccd1 vccd1 _19861_/X sky130_fd_sc_hd__clkbuf_1
X_18812_ _19555_/A _18812_/B vssd1 vssd1 vccd1 vccd1 _18812_/X sky130_fd_sc_hd__or2_1
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19792_ _19780_/X _19781_/X _19782_/X _19783_/X _19784_/X _19785_/X vssd1 vssd1 vccd1
+ vccd1 _19793_/A sky130_fd_sc_hd__mux4_1
XFILLER_122_496 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18743_ _18743_/A vssd1 vssd1 vccd1 vccd1 _26032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15955_ _15955_/A vssd1 vssd1 vccd1 vccd1 _15955_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14906_ _14906_/A vssd1 vssd1 vccd1 vccd1 _26481_/D sky130_fd_sc_hd__clkbuf_1
X_18674_ _26002_/Q _17753_/X _18674_/S vssd1 vssd1 vccd1 vccd1 _18675_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ _15887_/A vssd1 vssd1 vccd1 vccd1 _15886_/Y sky130_fd_sc_hd__inv_2
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _17671_/S vssd1 vssd1 vccd1 vccd1 _17634_/S sky130_fd_sc_hd__clkbuf_2
X_14837_ _14883_/S vssd1 vssd1 vccd1 vccd1 _14846_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_64_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17556_ _17460_/X _25854_/Q _17562_/S vssd1 vssd1 vccd1 vccd1 _17557_/A sky130_fd_sc_hd__mux2_1
X_14768_ _14768_/A vssd1 vssd1 vccd1 vccd1 _26536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16507_ _16815_/B _16545_/B vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__xor2_1
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13719_ _13900_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13719_/Y sky130_fd_sc_hd__nor2_1
X_17487_ _17487_/A vssd1 vssd1 vccd1 vccd1 _25830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14699_ _15771_/A _14699_/B vssd1 vssd1 vccd1 vccd1 _14699_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19226_ _19250_/A _19226_/B vssd1 vssd1 vccd1 vccd1 _19226_/X sky130_fd_sc_hd__or2_1
X_16438_ _16728_/A vssd1 vssd1 vccd1 vccd1 _16767_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19157_ _19250_/A _19157_/B vssd1 vssd1 vccd1 vccd1 _19157_/X sky130_fd_sc_hd__or2_1
XFILLER_145_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16369_ _16369_/A vssd1 vssd1 vccd1 vccd1 _16369_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18108_ _18108_/A _17978_/X vssd1 vssd1 vccd1 vccd1 _18108_/X sky130_fd_sc_hd__or2b_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19088_ _26692_/Q _26660_/Q _26628_/Q _26596_/Q _19015_/X _19087_/X vssd1 vssd1 vccd1
+ vccd1 _19088_/X sky130_fd_sc_hd__mux4_2
XFILLER_173_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18039_ _17888_/X _18035_/X _18038_/X _17894_/X vssd1 vssd1 vccd1 vccd1 _18039_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_536 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21050_ _21050_/A vssd1 vssd1 vccd1 vccd1 _21050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20001_ _20001_/A vssd1 vssd1 vccd1 vccd1 _20001_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21952_ _22000_/A vssd1 vssd1 vccd1 vccd1 _21952_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24740_ _24740_/A _24970_/A vssd1 vssd1 vccd1 vccd1 _24740_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ _20886_/X _20888_/X _20890_/X _20892_/X _20893_/X _20894_/X vssd1 vssd1 vccd1
+ vccd1 _20904_/A sky130_fd_sc_hd__mux4_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24671_ _27171_/Q _24671_/B vssd1 vssd1 vccd1 vccd1 _24671_/X sky130_fd_sc_hd__or2_1
X_21883_ _21899_/A vssd1 vssd1 vccd1 vccd1 _21883_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26410_ _20745_/X _26410_/D vssd1 vssd1 vccd1 vccd1 _26410_/Q sky130_fd_sc_hd__dfxtp_1
X_23622_ _23622_/A vssd1 vssd1 vccd1 vccd1 _27225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20834_ _20866_/A vssd1 vssd1 vccd1 vccd1 _20834_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27390_ _27394_/CLK _27390_/D vssd1 vssd1 vccd1 vccd1 _27390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26341_ _20505_/X _26341_/D vssd1 vssd1 vccd1 vccd1 _26341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23553_ _24877_/A _27207_/Q _23559_/S vssd1 vssd1 vccd1 vccd1 _23554_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20765_ _20765_/A vssd1 vssd1 vccd1 vccd1 _20765_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22504_ _22520_/A vssd1 vssd1 vccd1 vccd1 _22504_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26272_ _20261_/X _26272_/D vssd1 vssd1 vccd1 vccd1 _26272_/Q sky130_fd_sc_hd__dfxtp_1
X_23484_ input25/X _23482_/X _23483_/X _23474_/X vssd1 vssd1 vccd1 vccd1 _27186_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20696_ _20684_/X _20685_/X _20686_/X _20687_/X _20689_/X _20691_/X vssd1 vssd1 vccd1
+ vccd1 _20697_/A sky130_fd_sc_hd__mux4_1
XFILLER_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25223_ _25308_/A vssd1 vssd1 vccd1 vccd1 _25223_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_28011_ _28011_/A _15972_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_195_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22435_ _22435_/A vssd1 vssd1 vccd1 vccd1 _22435_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1077 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25154_ _27525_/Q _27493_/Q vssd1 vssd1 vccd1 vccd1 _25164_/A sky130_fd_sc_hd__nor2_1
X_22366_ _22433_/A vssd1 vssd1 vccd1 vccd1 _22366_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_544 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24105_ _24105_/A vssd1 vssd1 vccd1 vccd1 _27327_/D sky130_fd_sc_hd__clkbuf_1
X_21317_ _21301_/X _21302_/X _21303_/X _21304_/X _21307_/X _21310_/X vssd1 vssd1 vccd1
+ vccd1 _21318_/A sky130_fd_sc_hd__mux4_1
XFILLER_191_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25085_ _27839_/Q _27143_/Q _25888_/Q _25856_/Q _25061_/X _24975_/X vssd1 vssd1 vccd1
+ vccd1 _25085_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22297_ _22280_/X _22282_/X _22284_/X _22286_/X _22287_/X _22288_/X vssd1 vssd1 vccd1
+ vccd1 _22298_/A sky130_fd_sc_hd__mux4_1
XFILLER_123_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24036_ _27856_/Q _27160_/Q _25905_/Q _25873_/Q _24014_/X _23749_/X vssd1 vssd1 vccd1
+ vccd1 _24036_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21248_ _21248_/A vssd1 vssd1 vccd1 vccd1 _21248_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21179_ _21211_/A vssd1 vssd1 vccd1 vccd1 _21179_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_25987_ _25987_/CLK _25987_/D vssd1 vssd1 vccd1 vccd1 _25987_/Q sky130_fd_sc_hd__dfxtp_1
X_15740_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15740_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27726_ _27726_/CLK _27726_/D vssd1 vssd1 vccd1 vccd1 _27726_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _27819_/Q _12952_/B vssd1 vssd1 vccd1 vccd1 _12953_/A sky130_fd_sc_hd__and2_1
XFILLER_19_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24938_ _24938_/A vssd1 vssd1 vccd1 vccd1 _24938_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27657_ _27658_/CLK _27657_/D vssd1 vssd1 vccd1 vccd1 _27657_/Q sky130_fd_sc_hd__dfxtp_1
X_15671_ _15671_/A vssd1 vssd1 vccd1 vccd1 _26149_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _14511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24869_ _24873_/B _24869_/B vssd1 vssd1 vccd1 vccd1 _24870_/B sky130_fd_sc_hd__or2_1
XFILLER_93_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _14791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _17291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17410_/A vssd1 vssd1 vccd1 vccd1 _23109_/A sky130_fd_sc_hd__clkbuf_1
X_26608_ _21440_/X _26608_/D vssd1 vssd1 vccd1 vccd1 _26608_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _15695_/A _15695_/B _15695_/C _15407_/A vssd1 vssd1 vccd1 vccd1 _14639_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA_243 _25641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 _26824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18390_ _26288_/Q _26256_/Q _26224_/Q _26192_/Q _18301_/X _18324_/X vssd1 vssd1 vccd1
+ vccd1 _18390_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27588_ _27589_/CLK _27588_/D vssd1 vssd1 vccd1 vccd1 _27588_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_265 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _25838_/Q _26037_/Q _17341_/S vssd1 vssd1 vccd1 vccd1 _17341_/X sky130_fd_sc_hd__mux2_1
XANTENNA_287 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14553_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_298 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26539_ _21194_/X _26539_/D vssd1 vssd1 vccd1 vccd1 _26539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13504_ _26955_/Q _13487_/X _13482_/X _13503_/Y vssd1 vssd1 vccd1 vccd1 _26955_/D
+ sky130_fd_sc_hd__a31o_1
X_17272_ _27087_/Q _27119_/Q _17295_/S vssd1 vssd1 vccd1 vccd1 _17272_/X sky130_fd_sc_hd__mux2_1
X_14484_ _26632_/Q _14478_/X _14474_/X _14483_/Y vssd1 vssd1 vccd1 vccd1 _26632_/D
+ sky130_fd_sc_hd__a31o_1
X_19011_ _19107_/A _19011_/B _19011_/C vssd1 vssd1 vccd1 vccd1 _19012_/A sky130_fd_sc_hd__and3_1
XFILLER_146_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16223_ _23033_/A _16235_/B vssd1 vssd1 vccd1 vccd1 _16223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13435_ _25733_/B vssd1 vssd1 vccd1 vccd1 _13435_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16154_ _16152_/Y _16119_/X _16121_/X _14452_/A _16153_/Y vssd1 vssd1 vccd1 vccd1
+ _24300_/A sky130_fd_sc_hd__o221a_1
X_13366_ _14756_/A vssd1 vssd1 vccd1 vccd1 _13366_/X sky130_fd_sc_hd__buf_2
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15105_ _15105_/A vssd1 vssd1 vccd1 vccd1 _26400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_181_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16085_ _16699_/A vssd1 vssd1 vccd1 vccd1 _16621_/A sky130_fd_sc_hd__clkbuf_2
X_13297_ _13297_/A vssd1 vssd1 vccd1 vccd1 _27012_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15036_ _15775_/A _15043_/B vssd1 vssd1 vccd1 vccd1 _15036_/Y sky130_fd_sc_hd__nor2_1
X_19913_ _19913_/A vssd1 vssd1 vccd1 vccd1 _19913_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19844_ _19831_/X _19833_/X _19835_/X _19837_/X _19838_/X _19839_/X vssd1 vssd1 vccd1
+ vccd1 _19845_/A sky130_fd_sc_hd__mux4_1
XFILLER_123_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19775_ _19775_/A vssd1 vssd1 vccd1 vccd1 _19775_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1140 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16987_ _17380_/S vssd1 vssd1 vccd1 vccd1 _17307_/A sky130_fd_sc_hd__buf_2
XFILLER_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_561 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18726_ _18748_/A vssd1 vssd1 vccd1 vccd1 _18735_/S sky130_fd_sc_hd__buf_2
XFILLER_114_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15938_ _15956_/A vssd1 vssd1 vccd1 vccd1 _15943_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18657_ _25994_/Q _17728_/X _18663_/S vssd1 vssd1 vccd1 vccd1 _18658_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15869_ input1/X vssd1 vssd1 vccd1 vccd1 _15894_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ _17431_/X _25877_/Q _17612_/S vssd1 vssd1 vccd1 vccd1 _17609_/A sky130_fd_sc_hd__mux2_1
XFILLER_184_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18588_ _25434_/A vssd1 vssd1 vccd1 vccd1 _25474_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _17539_/A vssd1 vssd1 vccd1 vccd1 _25846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20550_ _20598_/A vssd1 vssd1 vccd1 vccd1 _20550_/X sky130_fd_sc_hd__clkbuf_1
X_19209_ _26953_/Q _26921_/Q _26889_/Q _26857_/Q _19208_/X _19116_/X vssd1 vssd1 vccd1
+ vccd1 _19209_/X sky130_fd_sc_hd__mux4_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater90 _25895_/CLK vssd1 vssd1 vccd1 vccd1 _27154_/CLK sky130_fd_sc_hd__clkbuf_1
X_20481_ _20513_/A vssd1 vssd1 vccd1 vccd1 _20481_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_28002__468 vssd1 vssd1 vccd1 vccd1 _28002__468/HI _28002_/A sky130_fd_sc_hd__conb_1
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22220_ _22220_/A vssd1 vssd1 vccd1 vccd1 _22220_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22151_ _22141_/X _22142_/X _22143_/X _22144_/X _22145_/X _22146_/X vssd1 vssd1 vccd1
+ vccd1 _22152_/A sky130_fd_sc_hd__mux4_1
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21102_ _21102_/A vssd1 vssd1 vccd1 vccd1 _21102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22082_ _22082_/A vssd1 vssd1 vccd1 vccd1 _22082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21033_ _21023_/X _21024_/X _21025_/X _21026_/X _21027_/X _21028_/X vssd1 vssd1 vccd1
+ vccd1 _21034_/A sky130_fd_sc_hd__mux4_1
X_25910_ _27266_/CLK _25910_/D vssd1 vssd1 vccd1 vccd1 _25910_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26890_ _22424_/X _26890_/D vssd1 vssd1 vccd1 vccd1 _26890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25841_ _26040_/CLK _25841_/D vssd1 vssd1 vccd1 vccd1 _25841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25772_ _25772_/A vssd1 vssd1 vccd1 vccd1 _27841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22984_ _22984_/A vssd1 vssd1 vccd1 vccd1 _22984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27511_ _27511_/CLK _27511_/D vssd1 vssd1 vccd1 vccd1 _27511_/Q sky130_fd_sc_hd__dfxtp_1
X_24723_ _27190_/Q _24725_/B vssd1 vssd1 vccd1 vccd1 _24723_/X sky130_fd_sc_hd__or2_1
XFILLER_28_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21935_ _22021_/A vssd1 vssd1 vccd1 vccd1 _22000_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_417 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27442_ _27442_/CLK _27442_/D vssd1 vssd1 vccd1 vccd1 _27442_/Q sky130_fd_sc_hd__dfxtp_1
X_21866_ _21914_/A vssd1 vssd1 vccd1 vccd1 _21866_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24654_ _27164_/Q _24658_/B vssd1 vssd1 vccd1 vccd1 _24654_/X sky130_fd_sc_hd__or2_1
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20817_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23605_ _23617_/A _23605_/B vssd1 vssd1 vccd1 vccd1 _23606_/A sky130_fd_sc_hd__and2_1
X_27373_ _27475_/CLK _27373_/D vssd1 vssd1 vccd1 vccd1 _27373_/Q sky130_fd_sc_hd__dfxtp_1
X_21797_ _21813_/A vssd1 vssd1 vccd1 vccd1 _21797_/X sky130_fd_sc_hd__clkbuf_2
X_24585_ _27653_/Q _24587_/B vssd1 vssd1 vccd1 vccd1 _24586_/A sky130_fd_sc_hd__and2_1
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26324_ _20443_/X _26324_/D vssd1 vssd1 vccd1 vccd1 _26324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20748_ _20738_/X _20739_/X _20740_/X _20741_/X _20742_/X _20743_/X vssd1 vssd1 vccd1
+ vccd1 _20749_/A sky130_fd_sc_hd__mux4_1
X_23536_ _27760_/Q _27202_/Q _23542_/S vssd1 vssd1 vccd1 vccd1 _23537_/B sky130_fd_sc_hd__mux2_1
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23467_ _27180_/Q _23470_/B vssd1 vssd1 vccd1 vccd1 _23467_/X sky130_fd_sc_hd__or2_1
X_26255_ _20207_/X _26255_/D vssd1 vssd1 vccd1 vccd1 _26255_/Q sky130_fd_sc_hd__dfxtp_1
X_20679_ _20679_/A vssd1 vssd1 vccd1 vccd1 _20679_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _27338_/Q _13193_/X _13194_/X _27306_/Q _13219_/X vssd1 vssd1 vccd1 vccd1
+ _16197_/A sky130_fd_sc_hd__a221o_1
X_22418_ _22434_/A vssd1 vssd1 vccd1 vccd1 _22418_/X sky130_fd_sc_hd__clkbuf_1
X_25206_ _25221_/A _25206_/B vssd1 vssd1 vccd1 vccd1 _25206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_195_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23398_ _24790_/A _27254_/Q _27245_/Q _24765_/A vssd1 vssd1 vccd1 vccd1 _23398_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_26186_ _19965_/X _26186_/D vssd1 vssd1 vccd1 vccd1 _26186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13151_ _27049_/Q _13150_/X _13167_/S vssd1 vssd1 vccd1 vccd1 _13152_/A sky130_fd_sc_hd__mux2_1
X_22349_ _22349_/A vssd1 vssd1 vccd1 vccd1 _22349_/X sky130_fd_sc_hd__clkbuf_1
X_25137_ _25129_/A _25126_/X _25129_/B _25127_/A vssd1 vssd1 vccd1 vccd1 _25138_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25068_ _25068_/A vssd1 vssd1 vccd1 vccd1 _27682_/D sky130_fd_sc_hd__clkbuf_1
X_13082_ _13082_/A vssd1 vssd1 vccd1 vccd1 _13082_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_877 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24019_ _24017_/X _24018_/X _24033_/S vssd1 vssd1 vccd1 vccd1 _24019_/X sky130_fd_sc_hd__mux2_1
X_16910_ _16662_/A _16662_/B _16550_/X vssd1 vssd1 vccd1 vccd1 _16911_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17890_ _18380_/A vssd1 vssd1 vccd1 vccd1 _17890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16841_ _16841_/A _16841_/B _16840_/X vssd1 vssd1 vccd1 vccd1 _16841_/X sky130_fd_sc_hd__or3b_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19560_ _19560_/A _19560_/B vssd1 vssd1 vccd1 vccd1 _19560_/X sky130_fd_sc_hd__or2_1
X_16772_ _16772_/A _16772_/B vssd1 vssd1 vccd1 vccd1 _16786_/A sky130_fd_sc_hd__xor2_1
X_13984_ _16289_/A vssd1 vssd1 vccd1 vccd1 _14359_/A sky130_fd_sc_hd__buf_2
XFILLER_20_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18511_ _18844_/A vssd1 vssd1 vccd1 vccd1 _18842_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15723_ _15723_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15723_/Y sky130_fd_sc_hd__nor2_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27709_ _27709_/CLK _27709_/D vssd1 vssd1 vccd1 vccd1 _27709_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12935_ _12935_/A vssd1 vssd1 vccd1 vccd1 _27858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19491_ _26549_/Q _26517_/Q _26485_/Q _27061_/Q _19401_/X _19445_/X vssd1 vssd1 vccd1
+ vccd1 _19491_/X sky130_fd_sc_hd__mux4_1
XFILLER_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18442_ _18440_/X _18441_/X _18488_/S vssd1 vssd1 vccd1 vccd1 _18442_/X sky130_fd_sc_hd__mux2_2
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15654_ _13133_/X _26156_/Q _15656_/S vssd1 vssd1 vccd1 vccd1 _15655_/A sky130_fd_sc_hd__mux2_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14605_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18373_ _17897_/X _18367_/X _18369_/X _18371_/X _18372_/X vssd1 vssd1 vccd1 vccd1
+ _18374_/C sky130_fd_sc_hd__a221o_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15585_/A vssd1 vssd1 vccd1 vccd1 _26187_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ _17324_/A vssd1 vssd1 vccd1 vccd1 _27941_/A sky130_fd_sc_hd__clkbuf_1
X_14536_ _14620_/B vssd1 vssd1 vccd1 vccd1 _14536_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17255_ _17216_/X _17255_/B vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__and2b_1
XFILLER_144_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14467_ _16277_/A vssd1 vssd1 vccd1 vccd1 _15736_/A sky130_fd_sc_hd__buf_2
XFILLER_179_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16206_ _16206_/A _16224_/B _16235_/C vssd1 vssd1 vccd1 vccd1 _16206_/X sky130_fd_sc_hd__and3_1
XFILLER_146_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13418_ _26971_/Q _13417_/X _13421_/S vssd1 vssd1 vccd1 vccd1 _13419_/A sky130_fd_sc_hd__mux2_1
XFILLER_190_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17186_ _27080_/Q _27112_/Q _17234_/S vssd1 vssd1 vccd1 vccd1 _17186_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14398_ _14398_/A vssd1 vssd1 vccd1 vccd1 _14398_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16137_ _16137_/A vssd1 vssd1 vccd1 vccd1 _16137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13349_ _13349_/A vssd1 vssd1 vccd1 vccd1 _26993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ _25975_/Q vssd1 vssd1 vccd1 vccd1 _16068_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15019_ _15756_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _15019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19827_ _19827_/A vssd1 vssd1 vccd1 vccd1 _19827_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19758_ _19745_/X _19747_/X _19749_/X _19751_/X _19752_/X _19753_/X vssd1 vssd1 vccd1
+ vccd1 _19759_/A sky130_fd_sc_hd__mux4_1
X_18709_ _26017_/Q _17699_/X _18713_/S vssd1 vssd1 vccd1 vccd1 _18710_/A sky130_fd_sc_hd__mux2_1
X_19689_ _19689_/A vssd1 vssd1 vccd1 vccd1 _19689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21720_ _21720_/A vssd1 vssd1 vccd1 vccd1 _21720_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_681 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21651_ _21651_/A vssd1 vssd1 vccd1 vccd1 _21725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20602_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20672_/A sky130_fd_sc_hd__buf_2
XFILLER_162_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24370_ _27567_/Q _24372_/B vssd1 vssd1 vccd1 vccd1 _24371_/A sky130_fd_sc_hd__and2_1
X_21582_ _21648_/A vssd1 vssd1 vccd1 vccd1 _21582_/X sky130_fd_sc_hd__clkbuf_1
X_23321_ _23321_/A _23321_/B _23321_/C _23321_/D vssd1 vssd1 vccd1 vccd1 _23322_/B
+ sky130_fd_sc_hd__or4_1
X_20533_ _20599_/A vssd1 vssd1 vccd1 vccd1 _20533_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26040_ _26040_/CLK _26040_/D vssd1 vssd1 vccd1 vccd1 _26040_/Q sky130_fd_sc_hd__dfxtp_1
X_23252_ _17523_/X _27161_/Q _23252_/S vssd1 vssd1 vccd1 vccd1 _23253_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_497 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20464_ _20512_/A vssd1 vssd1 vccd1 vccd1 _20464_/X sky130_fd_sc_hd__clkbuf_1
X_22203_ _22194_/X _22196_/X _22198_/X _22200_/X _22201_/X _22202_/X vssd1 vssd1 vccd1
+ vccd1 _22204_/A sky130_fd_sc_hd__mux4_1
XFILLER_118_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23183_ _23239_/A vssd1 vssd1 vccd1 vccd1 _23252_/S sky130_fd_sc_hd__buf_2
XFILLER_133_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20395_ _20427_/A vssd1 vssd1 vccd1 vccd1 _20395_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22134_ _22134_/A vssd1 vssd1 vccd1 vccd1 _22134_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27991_ _27991_/A _15891_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_88_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_517 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22065_ _22051_/X _22052_/X _22053_/X _22054_/X _22055_/X _22056_/X vssd1 vssd1 vccd1
+ vccd1 _22066_/A sky130_fd_sc_hd__mux4_1
X_26942_ _22604_/X _26942_/D vssd1 vssd1 vccd1 vccd1 _26942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21016_ _21016_/A vssd1 vssd1 vccd1 vccd1 _21016_/X sky130_fd_sc_hd__clkbuf_1
X_26873_ _22362_/X _26873_/D vssd1 vssd1 vccd1 vccd1 _26873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25824_ _25991_/CLK _25824_/D vssd1 vssd1 vccd1 vccd1 _25824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_637 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25755_ _17450_/X _27834_/Q _25757_/S vssd1 vssd1 vccd1 vccd1 _25756_/A sky130_fd_sc_hd__mux2_1
X_22967_ _22955_/X _22956_/X _22957_/X _22958_/X _22960_/X _22962_/X vssd1 vssd1 vccd1
+ vccd1 _22968_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24706_ _24400_/A _24700_/X _24705_/X _24703_/X vssd1 vssd1 vccd1 vccd1 _27599_/D
+ sky130_fd_sc_hd__o211a_1
X_21918_ _21986_/A vssd1 vssd1 vccd1 vccd1 _21918_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_188_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25686_ _25686_/A vssd1 vssd1 vccd1 vccd1 _25686_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22898_ _22898_/A vssd1 vssd1 vccd1 vccd1 _22898_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27425_ _27425_/CLK _27425_/D vssd1 vssd1 vccd1 vccd1 _27425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24637_ _24637_/A vssd1 vssd1 vccd1 vccd1 _27576_/D sky130_fd_sc_hd__clkbuf_1
X_21849_ _22021_/A vssd1 vssd1 vccd1 vccd1 _21914_/A sky130_fd_sc_hd__buf_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15370_ _15392_/A vssd1 vssd1 vccd1 vccd1 _15379_/S sky130_fd_sc_hd__clkbuf_2
X_27356_ _27356_/CLK _27356_/D vssd1 vssd1 vccd1 vccd1 _27356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24568_ _27645_/Q _24576_/B vssd1 vssd1 vccd1 vccd1 _24569_/A sky130_fd_sc_hd__and2_1
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14321_ _26684_/Q _14310_/X _14311_/X _14320_/Y vssd1 vssd1 vccd1 vccd1 _26684_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26307_ _20387_/X _26307_/D vssd1 vssd1 vccd1 vccd1 _26307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23519_ _23519_/A vssd1 vssd1 vccd1 vccd1 _27197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27287_ _27423_/CLK _27287_/D vssd1 vssd1 vccd1 vccd1 _27287_/Q sky130_fd_sc_hd__dfxtp_1
X_24499_ _24638_/A vssd1 vssd1 vccd1 vccd1 _24499_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17040_ _27829_/Q _27133_/Q _25878_/Q _25846_/Q _17015_/X _16989_/X vssd1 vssd1 vccd1
+ vccd1 _17040_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14252_ _14340_/A _14263_/B vssd1 vssd1 vccd1 vccd1 _14252_/Y sky130_fd_sc_hd__nor2_1
X_26238_ _20143_/X _26238_/D vssd1 vssd1 vccd1 vccd1 _26238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13203_ _16212_/A vssd1 vssd1 vccd1 vccd1 _14791_/A sky130_fd_sc_hd__buf_2
X_14183_ _26735_/Q _14173_/X _14181_/X _14182_/Y vssd1 vssd1 vccd1 vccd1 _26735_/D
+ sky130_fd_sc_hd__a31o_1
X_26169_ _19897_/X _26169_/D vssd1 vssd1 vccd1 vccd1 _26169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_641 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13134_ _27052_/Q _13133_/X _13140_/S vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__mux2_1
X_18991_ _24511_/A vssd1 vssd1 vccd1 vccd1 _19473_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _27300_/Q _13125_/B vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__and2_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17942_ _26525_/Q _26493_/Q _26461_/Q _27037_/Q _17841_/X _17843_/X vssd1 vssd1 vccd1
+ vccd1 _17942_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater208 _27417_/CLK vssd1 vssd1 vccd1 vccd1 _25987_/CLK sky130_fd_sc_hd__clkbuf_1
X_17873_ _18358_/A vssd1 vssd1 vccd1 vccd1 _17873_/X sky130_fd_sc_hd__buf_2
Xrepeater219 _27398_/CLK vssd1 vssd1 vccd1 vccd1 _27397_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_572 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16824_ _16824_/A _16824_/B vssd1 vssd1 vccd1 vccd1 _16824_/Y sky130_fd_sc_hd__nand2_1
X_19612_ _19612_/A vssd1 vssd1 vccd1 vccd1 _19612_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19543_ _26296_/Q _26264_/Q _26232_/Q _26200_/Q _18908_/X _19486_/X vssd1 vssd1 vccd1
+ vccd1 _19543_/X sky130_fd_sc_hd__mux4_1
XFILLER_111_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16755_ _16755_/A _16756_/B vssd1 vssd1 vccd1 vccd1 _16755_/Y sky130_fd_sc_hd__nand2_1
X_13967_ _14346_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _13967_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15706_ _15712_/A vssd1 vssd1 vccd1 vccd1 _15761_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19474_ _26837_/Q _26805_/Q _26773_/Q _26741_/Q _18788_/X _19407_/X vssd1 vssd1 vccd1
+ vccd1 _19475_/B sky130_fd_sc_hd__mux4_1
X_16686_ _16686_/A _16686_/B vssd1 vssd1 vccd1 vccd1 _16686_/Y sky130_fd_sc_hd__nand2_1
X_13898_ _26827_/Q _13893_/X _13886_/X _13897_/Y vssd1 vssd1 vccd1 vccd1 _26827_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18425_ _18425_/A vssd1 vssd1 vccd1 vccd1 _18425_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ _13086_/X _26164_/Q _15645_/S vssd1 vssd1 vccd1 vccd1 _15638_/A sky130_fd_sc_hd__mux2_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18356_ _26959_/Q _26927_/Q _26895_/Q _26863_/Q _18244_/X _18269_/X vssd1 vssd1 vccd1
+ vccd1 _18356_/X sky130_fd_sc_hd__mux4_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _15568_/A vssd1 vssd1 vccd1 vccd1 _26195_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17307_ _17307_/A vssd1 vssd1 vccd1 vccd1 _17355_/S sky130_fd_sc_hd__clkbuf_2
X_14519_ _15771_/A _14519_/B vssd1 vssd1 vccd1 vccd1 _14519_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18287_ _18398_/A _18287_/B _18287_/C vssd1 vssd1 vccd1 vccd1 _18288_/A sky130_fd_sc_hd__and3_1
XFILLER_174_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15499_ _13105_/X _26225_/Q _15501_/S vssd1 vssd1 vccd1 vccd1 _15500_/A sky130_fd_sc_hd__mux2_1
X_17238_ _17299_/A vssd1 vssd1 vccd1 vccd1 _17238_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17169_ _17380_/S vssd1 vssd1 vccd1 vccd1 _17219_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20180_ _20266_/A vssd1 vssd1 vccd1 vccd1 _20248_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23870_ _23868_/X _23869_/X _23893_/S vssd1 vssd1 vccd1 vccd1 _23870_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22821_ _22869_/A vssd1 vssd1 vccd1 vccd1 _22821_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25540_ _25540_/A vssd1 vssd1 vccd1 vccd1 _25540_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22752_ _22784_/A vssd1 vssd1 vccd1 vccd1 _22752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_837 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21703_ _21689_/X _21690_/X _21691_/X _21692_/X _21693_/X _21694_/X vssd1 vssd1 vccd1
+ vccd1 _21704_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22683_ _22699_/A vssd1 vssd1 vccd1 vccd1 _22683_/X sky130_fd_sc_hd__clkbuf_1
X_25471_ _25456_/X _25461_/X _25462_/X _24849_/B _25463_/X vssd1 vssd1 vccd1 vccd1
+ _25471_/X sky130_fd_sc_hd__o311a_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28008__474 vssd1 vssd1 vccd1 vccd1 _28008__474/HI _28008_/A sky130_fd_sc_hd__conb_1
X_27210_ _27856_/CLK _27210_/D vssd1 vssd1 vccd1 vccd1 _27210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21634_ _21650_/A vssd1 vssd1 vccd1 vccd1 _21634_/X sky130_fd_sc_hd__clkbuf_1
X_24422_ _27611_/Q _24422_/B vssd1 vssd1 vccd1 vccd1 _24423_/A sky130_fd_sc_hd__and2_1
XFILLER_100_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27141_ _27141_/CLK _27141_/D vssd1 vssd1 vccd1 vccd1 _27141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21565_ _21651_/A vssd1 vssd1 vccd1 vccd1 _21635_/A sky130_fd_sc_hd__clkbuf_2
X_24353_ _27559_/Q _24361_/B vssd1 vssd1 vccd1 vccd1 _24354_/A sky130_fd_sc_hd__and2_1
XFILLER_21_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23304_ _27734_/Q _23267_/Y _27749_/Q _23301_/Y _23303_/Y vssd1 vssd1 vccd1 vccd1
+ _23309_/B sky130_fd_sc_hd__a221o_1
X_20516_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20586_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24284_ _24284_/A _24287_/B vssd1 vssd1 vccd1 vccd1 _24285_/A sky130_fd_sc_hd__and2_1
X_27072_ _27105_/CLK _27072_/D vssd1 vssd1 vccd1 vccd1 _27072_/Q sky130_fd_sc_hd__dfxtp_1
X_21496_ _21562_/A vssd1 vssd1 vccd1 vccd1 _21496_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1068 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23235_ _17498_/X _27153_/Q _23237_/S vssd1 vssd1 vccd1 vccd1 _23236_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26023_ _27112_/CLK _26023_/D vssd1 vssd1 vccd1 vccd1 _26023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20447_ _20513_/A vssd1 vssd1 vccd1 vccd1 _20447_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23166_ _23166_/A vssd1 vssd1 vccd1 vccd1 _27122_/D sky130_fd_sc_hd__clkbuf_1
X_20378_ _20426_/A vssd1 vssd1 vccd1 vccd1 _20378_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22117_ _22103_/X _22106_/X _22109_/X _22112_/X _22113_/X _22114_/X vssd1 vssd1 vccd1
+ vccd1 _22118_/A sky130_fd_sc_hd__mux4_1
XFILLER_0_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23097_ _27092_/Q _17760_/X _23103_/S vssd1 vssd1 vccd1 vccd1 _23098_/A sky130_fd_sc_hd__mux2_1
X_27974_ _27974_/A _15936_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
XFILLER_125_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22048_ _22048_/A vssd1 vssd1 vccd1 vccd1 _22048_/X sky130_fd_sc_hd__clkbuf_1
X_26925_ _22552_/X _26925_/D vssd1 vssd1 vccd1 vccd1 _26925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26856_ _22308_/X _26856_/D vssd1 vssd1 vccd1 vccd1 _26856_/Q sky130_fd_sc_hd__dfxtp_1
X_14870_ _14870_/A vssd1 vssd1 vccd1 vccd1 _14879_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_47_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13821_ _13913_/A _13825_/B vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__nor2_1
X_25807_ _25721_/X _25722_/X _25723_/X _25724_/X _25725_/X _25726_/X vssd1 vssd1 vccd1
+ vccd1 _25808_/A sky130_fd_sc_hd__mux4_2
X_26787_ _22062_/X _26787_/D vssd1 vssd1 vccd1 vccd1 _26787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23999_ _27788_/Q vssd1 vssd1 vccd1 vccd1 _24033_/S sky130_fd_sc_hd__clkbuf_2
X_16540_ _16802_/A _16540_/B vssd1 vssd1 vccd1 vccd1 _16616_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13752_ _26878_/Q _13750_/X _13745_/X _13751_/Y vssd1 vssd1 vccd1 vccd1 _26878_/D
+ sky130_fd_sc_hd__a31o_1
X_25738_ _17408_/X _27826_/Q _25746_/S vssd1 vssd1 vccd1 vccd1 _25739_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16471_ _16778_/B _16471_/B vssd1 vssd1 vccd1 vccd1 _16609_/A sky130_fd_sc_hd__or2_1
XFILLER_189_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13683_ _13861_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13683_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25669_ _25654_/X _25656_/X _25658_/X _25660_/X _25661_/X _25662_/X vssd1 vssd1 vccd1
+ vccd1 _25670_/A sky130_fd_sc_hd__mux4_1
X_18210_ _26280_/Q _26248_/Q _26216_/Q _26184_/Q _18185_/X _18209_/X vssd1 vssd1 vccd1
+ vccd1 _18210_/X sky130_fd_sc_hd__mux4_1
X_15422_ _15422_/A vssd1 vssd1 vccd1 vccd1 _26260_/D sky130_fd_sc_hd__clkbuf_1
X_27408_ _27408_/CLK _27408_/D vssd1 vssd1 vccd1 vccd1 _27408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19190_ _19261_/A _19190_/B vssd1 vssd1 vccd1 vccd1 _19190_/X sky130_fd_sc_hd__or2_1
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18141_ _18141_/A vssd1 vssd1 vccd1 vccd1 _18141_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _14734_/X _26290_/Q _15357_/S vssd1 vssd1 vccd1 vccd1 _15354_/A sky130_fd_sc_hd__mux2_1
X_27339_ _27341_/CLK _27339_/D vssd1 vssd1 vccd1 vccd1 _27339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ _14304_/A vssd1 vssd1 vccd1 vccd1 _14316_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18072_ _26530_/Q _26498_/Q _26466_/Q _27042_/Q _17964_/X _17986_/X vssd1 vssd1 vccd1
+ vccd1 _18072_/X sky130_fd_sc_hd__mux4_1
X_15284_ _26320_/Q _13350_/X _15284_/S vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__mux2_1
X_17023_ _16985_/X _17016_/X _17020_/X _17022_/X vssd1 vssd1 vccd1 vccd1 _17023_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_172_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14235_ _26714_/Q _14225_/X _14158_/B _14234_/Y vssd1 vssd1 vccd1 vccd1 _26714_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14166_ _14166_/A vssd1 vssd1 vccd1 vccd1 _14220_/A sky130_fd_sc_hd__buf_2
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13241_/S vssd1 vssd1 vccd1 vccd1 _13140_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _26766_/Q _14090_/X _14093_/X _14096_/Y vssd1 vssd1 vccd1 vccd1 _26766_/D
+ sky130_fd_sc_hd__a31o_1
X_18974_ _19465_/A vssd1 vssd1 vccd1 vccd1 _18974_/X sky130_fd_sc_hd__buf_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17925_ _18437_/A vssd1 vssd1 vccd1 vccd1 _18056_/S sky130_fd_sc_hd__clkbuf_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13048_ _15551_/A vssd1 vssd1 vccd1 vccd1 _15695_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17856_ _18238_/A vssd1 vssd1 vccd1 vccd1 _17856_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16807_ _16807_/A _16807_/B vssd1 vssd1 vccd1 vccd1 _16807_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17787_ _27593_/Q vssd1 vssd1 vccd1 vccd1 _17898_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14999_ _15738_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _14999_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16738_ _16738_/A _16738_/B vssd1 vssd1 vccd1 vccd1 _16738_/Y sky130_fd_sc_hd__nand2_1
X_19526_ _19485_/X _19525_/X _19488_/X vssd1 vssd1 vccd1 vccd1 _19526_/X sky130_fd_sc_hd__o21a_1
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19457_ _27819_/Q _26580_/Q _26452_/Q _26132_/Q _19414_/X _18831_/X vssd1 vssd1 vccd1
+ vccd1 _19457_/X sky130_fd_sc_hd__mux4_1
X_16669_ _16077_/A _16670_/A _16809_/B _16650_/A vssd1 vssd1 vccd1 vccd1 _16669_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_179_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18408_ _18408_/A vssd1 vssd1 vccd1 vccd1 _18408_/X sky130_fd_sc_hd__clkbuf_2
X_19388_ _19273_/X _19386_/X _19387_/X vssd1 vssd1 vccd1 vccd1 _19388_/X sky130_fd_sc_hd__o21a_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18339_ _27813_/Q _26574_/Q _26446_/Q _26126_/Q _18011_/A _18427_/A vssd1 vssd1 vccd1
+ vccd1 _18339_/X sky130_fd_sc_hd__mux4_2
XFILLER_175_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21350_ _21350_/A vssd1 vssd1 vccd1 vccd1 _21350_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20301_ _20301_/A vssd1 vssd1 vccd1 vccd1 _20301_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21281_ _21269_/X _21270_/X _21271_/X _21272_/X _21273_/X _21274_/X vssd1 vssd1 vccd1
+ vccd1 _21282_/A sky130_fd_sc_hd__mux4_1
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23020_ _23020_/A vssd1 vssd1 vccd1 vccd1 _23020_/X sky130_fd_sc_hd__clkbuf_1
X_20232_ _20248_/A vssd1 vssd1 vccd1 vccd1 _20232_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20163_ _20163_/A vssd1 vssd1 vccd1 vccd1 _20163_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20094_ _20266_/A vssd1 vssd1 vccd1 vccd1 _20162_/A sky130_fd_sc_hd__buf_2
X_24971_ _27671_/Q _24838_/A _24970_/Y _24663_/A vssd1 vssd1 vccd1 vccd1 _27671_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26710_ _21800_/X _26710_/D vssd1 vssd1 vccd1 vccd1 _26710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23922_ _25929_/Q _25995_/Q _25828_/Q _26027_/Q _23899_/X _23882_/X vssd1 vssd1 vccd1
+ vccd1 _23922_/X sky130_fd_sc_hd__mux4_1
X_27690_ _27690_/CLK _27690_/D vssd1 vssd1 vccd1 vccd1 _27690_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26641_ _21554_/X _26641_/D vssd1 vssd1 vccd1 vccd1 _26641_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23853_ _25922_/Q _25988_/Q _25821_/Q _26020_/Q _23852_/X _23835_/X vssd1 vssd1 vccd1
+ vccd1 _23853_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22804_ _22870_/A vssd1 vssd1 vccd1 vccd1 _22804_/X sky130_fd_sc_hd__clkbuf_1
X_26572_ _21316_/X _26572_/D vssd1 vssd1 vccd1 vccd1 _26572_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _21028_/A vssd1 vssd1 vccd1 vccd1 _20996_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_23784_ _23740_/X _23782_/X _23783_/X _23768_/X vssd1 vssd1 vccd1 vccd1 _27273_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25523_ _25553_/A vssd1 vssd1 vccd1 vccd1 _25523_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22735_ _22783_/A vssd1 vssd1 vccd1 vccd1 _22735_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_492 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25454_ _24737_/A _25431_/X _25450_/Y _25453_/X _25446_/X vssd1 vssd1 vccd1 vccd1
+ _27756_/D sky130_fd_sc_hd__a221oi_1
X_22666_ _22698_/A vssd1 vssd1 vccd1 vccd1 _22666_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24405_ _24405_/A _24411_/B vssd1 vssd1 vccd1 vccd1 _24406_/A sky130_fd_sc_hd__and2_1
XFILLER_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21617_ _21649_/A vssd1 vssd1 vccd1 vccd1 _21617_/X sky130_fd_sc_hd__clkbuf_1
X_25385_ _27732_/Q input43/X _25391_/S vssd1 vssd1 vccd1 vccd1 _25386_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22597_ _22597_/A vssd1 vssd1 vccd1 vccd1 _22597_/X sky130_fd_sc_hd__clkbuf_2
X_27124_ _27124_/CLK _27124_/D vssd1 vssd1 vccd1 vccd1 _27124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24336_ _24336_/A vssd1 vssd1 vccd1 vccd1 _27451_/D sky130_fd_sc_hd__clkbuf_1
X_21548_ _21564_/A vssd1 vssd1 vccd1 vccd1 _21548_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27055_ _23000_/X _27055_/D vssd1 vssd1 vccd1 vccd1 _27055_/Q sky130_fd_sc_hd__dfxtp_1
X_21479_ _21651_/A vssd1 vssd1 vccd1 vccd1 _21549_/A sky130_fd_sc_hd__clkbuf_2
X_24267_ _24267_/A _24287_/B vssd1 vssd1 vccd1 vccd1 _24268_/A sky130_fd_sc_hd__and2_1
XFILLER_181_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14020_ _14493_/A vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__buf_2
X_26006_ _26007_/CLK _26006_/D vssd1 vssd1 vccd1 vccd1 _26006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23218_ _17472_/X _27145_/Q _23226_/S vssd1 vssd1 vccd1 vccd1 _23219_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24198_ _24238_/A vssd1 vssd1 vccd1 vccd1 _24363_/A sky130_fd_sc_hd__buf_2
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23149_ _23149_/A vssd1 vssd1 vccd1 vccd1 _27114_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_953 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27957_ _27957_/A _15920_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
X_15971_ _15973_/A vssd1 vssd1 vccd1 vccd1 _15971_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17710_ _25922_/Q _17708_/X _17722_/S vssd1 vssd1 vccd1 vccd1 _17711_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26908_ _22484_/X _26908_/D vssd1 vssd1 vccd1 vccd1 _26908_/Q sky130_fd_sc_hd__dfxtp_1
X_14922_ _14922_/A vssd1 vssd1 vccd1 vccd1 _26474_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18690_ _18690_/A vssd1 vssd1 vccd1 vccd1 _26009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17641_ _17479_/X _25892_/Q _17645_/S vssd1 vssd1 vccd1 vccd1 _17642_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26839_ _22244_/X _26839_/D vssd1 vssd1 vccd1 vccd1 _26839_/Q sky130_fd_sc_hd__dfxtp_1
X_14853_ _26504_/Q _13376_/X _14857_/S vssd1 vssd1 vccd1 vccd1 _14854_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ _13897_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17572_ _17572_/A vssd1 vssd1 vccd1 vccd1 _25861_/D sky130_fd_sc_hd__clkbuf_1
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _26531_/D sky130_fd_sc_hd__clkbuf_1
X_19311_ _27602_/Q vssd1 vssd1 vccd1 vccd1 _19312_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_16523_ _16826_/A vssd1 vssd1 vccd1 vccd1 _16908_/A sky130_fd_sc_hd__inv_2
X_13735_ _13915_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13735_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19242_ _19401_/A vssd1 vssd1 vccd1 vccd1 _19242_/X sky130_fd_sc_hd__buf_2
XFILLER_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16454_ _16422_/A _16256_/B _16256_/C _16459_/A _16360_/A vssd1 vssd1 vccd1 vccd1
+ _16455_/B sky130_fd_sc_hd__o41a_1
X_13666_ _13936_/A _13670_/B vssd1 vssd1 vccd1 vccd1 _13666_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15405_ _14810_/X _26266_/Q _15405_/S vssd1 vssd1 vccd1 vccd1 _15406_/A sky130_fd_sc_hd__mux2_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19173_ _19171_/X _19172_/X _19173_/S vssd1 vssd1 vccd1 vccd1 _19173_/X sky130_fd_sc_hd__mux2_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _17420_/B _16490_/B vssd1 vssd1 vccd1 vccd1 _16385_/Y sky130_fd_sc_hd__nor2_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _13868_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13597_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18124_ _18146_/A _18124_/B _18124_/C vssd1 vssd1 vccd1 vccd1 _18125_/A sky130_fd_sc_hd__and3_1
XFILLER_145_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15336_ _15392_/A vssd1 vssd1 vccd1 vccd1 _15405_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_157_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18055_ _26946_/Q _26914_/Q _26882_/Q _26850_/Q _17922_/X _17951_/X vssd1 vssd1 vccd1
+ vccd1 _18055_/X sky130_fd_sc_hd__mux4_2
X_15267_ _26328_/Q _13325_/X _15273_/S vssd1 vssd1 vccd1 vccd1 _15268_/A sky130_fd_sc_hd__mux2_1
XANTENNA_2 _20577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17006_ input38/X vssd1 vssd1 vccd1 vccd1 _17048_/S sky130_fd_sc_hd__clkbuf_2
X_14218_ _14396_/A _14226_/B vssd1 vssd1 vccd1 vccd1 _14218_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_461 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15198_ _15198_/A vssd1 vssd1 vccd1 vccd1 _26359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ _15695_/D _14149_/B vssd1 vssd1 vccd1 vccd1 _14166_/A sky130_fd_sc_hd__or2_1
XFILLER_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18957_ _27601_/Q vssd1 vssd1 vccd1 vccd1 _19488_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17908_ _17959_/A vssd1 vssd1 vccd1 vccd1 _24386_/A sky130_fd_sc_hd__clkbuf_4
X_18888_ _26396_/Q _26364_/Q _26332_/Q _26300_/Q _18887_/X _18826_/X vssd1 vssd1 vccd1
+ vccd1 _18888_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17839_ _17830_/X _17836_/X _17838_/X vssd1 vssd1 vccd1 vccd1 _17839_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20850_ _20866_/A vssd1 vssd1 vccd1 vccd1 _20850_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19509_ _26422_/Q _26390_/Q _26358_/Q _26326_/Q _19465_/X _18795_/X vssd1 vssd1 vccd1
+ vccd1 _19509_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20781_ _20781_/A vssd1 vssd1 vccd1 vccd1 _20781_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22520_ _22520_/A vssd1 vssd1 vccd1 vccd1 _22520_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22451_ _22451_/A vssd1 vssd1 vccd1 vccd1 _22519_/A sky130_fd_sc_hd__buf_2
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_687 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21402_ _21402_/A vssd1 vssd1 vccd1 vccd1 _21402_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22382_ _22382_/A vssd1 vssd1 vccd1 vccd1 _22382_/X sky130_fd_sc_hd__clkbuf_1
X_25170_ _25170_/A _25169_/Y vssd1 vssd1 vccd1 vccd1 _25173_/A sky130_fd_sc_hd__or2b_1
XFILLER_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21333_ _21322_/X _21324_/X _21326_/X _21328_/X _21329_/X _21330_/X vssd1 vssd1 vccd1
+ vccd1 _21334_/A sky130_fd_sc_hd__mux4_1
X_24121_ _24121_/A vssd1 vssd1 vccd1 vccd1 _27334_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1185 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21264_ _21264_/A vssd1 vssd1 vccd1 vccd1 _21264_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24052_ _24063_/A vssd1 vssd1 vccd1 vccd1 _24061_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20215_ _20215_/A vssd1 vssd1 vccd1 vccd1 _20215_/X sky130_fd_sc_hd__clkbuf_1
X_23003_ _22993_/X _22994_/X _22995_/X _22996_/X _22997_/X _22998_/X vssd1 vssd1 vccd1
+ vccd1 _23004_/A sky130_fd_sc_hd__mux4_1
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21195_ _21211_/A vssd1 vssd1 vccd1 vccd1 _21195_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27811_ _25688_/X _27811_/D vssd1 vssd1 vccd1 vccd1 _27811_/Q sky130_fd_sc_hd__dfxtp_1
X_20146_ _20162_/A vssd1 vssd1 vccd1 vccd1 _20146_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27742_ _27745_/CLK _27742_/D vssd1 vssd1 vccd1 vccd1 _27742_/Q sky130_fd_sc_hd__dfxtp_1
X_20077_ _20077_/A vssd1 vssd1 vccd1 vccd1 _20077_/X sky130_fd_sc_hd__clkbuf_1
X_24954_ _25601_/A _24954_/B _24954_/C vssd1 vssd1 vccd1 vccd1 _24960_/B sky130_fd_sc_hd__and3_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23905_ _27788_/Q vssd1 vssd1 vccd1 vccd1 _23940_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27673_ _27678_/CLK _27673_/D vssd1 vssd1 vccd1 vccd1 _27964_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24885_ _24935_/A vssd1 vssd1 vccd1 vccd1 _24885_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater380 _27563_/CLK vssd1 vssd1 vccd1 vccd1 _27225_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26624_ _21492_/X _26624_/D vssd1 vssd1 vccd1 vccd1 _26624_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater391 _27447_/CLK vssd1 vssd1 vccd1 vccd1 _27222_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_73_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23836_ _25920_/Q _25986_/Q _25819_/Q _26018_/Q _23804_/X _23835_/X vssd1 vssd1 vccd1
+ vccd1 _23836_/X sky130_fd_sc_hd__mux4_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26555_ _21260_/X _26555_/D vssd1 vssd1 vccd1 vccd1 _26555_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23767_ _24063_/A vssd1 vssd1 vccd1 vccd1 _23864_/A sky130_fd_sc_hd__buf_2
X_20979_ _21027_/A vssd1 vssd1 vccd1 vccd1 _20979_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13520_ _16243_/A vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__clkbuf_2
X_25506_ _25487_/X _25492_/X _25493_/X _24878_/B _25494_/X vssd1 vssd1 vccd1 vccd1
+ _25506_/X sky130_fd_sc_hd__o311a_1
XFILLER_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22718_ _22784_/A vssd1 vssd1 vccd1 vccd1 _22718_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_186_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26486_ _21016_/X _26486_/D vssd1 vssd1 vccd1 vccd1 _26486_/Q sky130_fd_sc_hd__dfxtp_1
X_23698_ _23698_/A vssd1 vssd1 vccd1 vccd1 _27253_/D sky130_fd_sc_hd__clkbuf_1
X_25437_ _25437_/A vssd1 vssd1 vccd1 vccd1 _25560_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13451_ _13530_/A vssd1 vssd1 vccd1 vccd1 _13451_/X sky130_fd_sc_hd__buf_4
X_22649_ _22697_/A vssd1 vssd1 vccd1 vccd1 _22649_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16170_ _27529_/Q _16034_/A vssd1 vssd1 vccd1 vccd1 _16170_/X sky130_fd_sc_hd__or2b_1
XFILLER_167_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13382_ _16240_/A vssd1 vssd1 vccd1 vccd1 _13382_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25368_ _25368_/A vssd1 vssd1 vccd1 vccd1 _27724_/D sky130_fd_sc_hd__clkbuf_1
X_27107_ _27413_/CLK _27107_/D vssd1 vssd1 vccd1 vccd1 _27107_/Q sky130_fd_sc_hd__dfxtp_1
X_15121_ _26393_/Q _13319_/X _15129_/S vssd1 vssd1 vccd1 vccd1 _15122_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24319_ _24330_/A vssd1 vssd1 vccd1 vccd1 _24328_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_127_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25299_ _25299_/A vssd1 vssd1 vccd1 vccd1 _25299_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27038_ _22936_/X _27038_/D vssd1 vssd1 vccd1 vccd1 _27038_/Q sky130_fd_sc_hd__dfxtp_1
X_15052_ _15052_/A vssd1 vssd1 vccd1 vccd1 _26424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14003_ _14372_/A _14010_/B vssd1 vssd1 vccd1 vccd1 _14003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19860_ _19850_/X _19851_/X _19852_/X _19853_/X _19854_/X _19855_/X vssd1 vssd1 vccd1
+ vccd1 _19861_/A sky130_fd_sc_hd__mux4_1
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18811_ _26138_/Q _26074_/Q _27002_/Q _26970_/Q _18807_/X _18810_/X vssd1 vssd1 vccd1
+ vccd1 _18812_/B sky130_fd_sc_hd__mux4_1
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19791_ _19791_/A vssd1 vssd1 vccd1 vccd1 _19791_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_795 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18742_ _26032_/Q _17747_/X _18746_/S vssd1 vssd1 vccd1 vccd1 _18743_/A sky130_fd_sc_hd__mux2_1
X_15954_ _15955_/A vssd1 vssd1 vccd1 vccd1 _15954_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14905_ _14737_/X _26481_/Q _14907_/S vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__mux2_1
X_18673_ _18673_/A vssd1 vssd1 vccd1 vccd1 _26001_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _15887_/A vssd1 vssd1 vccd1 vccd1 _15885_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ _14836_/A vssd1 vssd1 vccd1 vccd1 _26512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17624_ _17624_/A vssd1 vssd1 vccd1 vccd1 _25884_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _17555_/A vssd1 vssd1 vccd1 vccd1 _25853_/D sky130_fd_sc_hd__clkbuf_1
X_14767_ _14766_/X _26536_/Q _14773_/S vssd1 vssd1 vccd1 vccd1 _14768_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16506_ _16633_/A _16506_/B vssd1 vssd1 vccd1 vccd1 _16545_/B sky130_fd_sc_hd__xnor2_1
X_13718_ _13745_/A vssd1 vssd1 vccd1 vccd1 _13718_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17486_ _17485_/X _25830_/Q _17486_/S vssd1 vssd1 vccd1 vccd1 _17487_/A sky130_fd_sc_hd__mux2_1
X_14698_ _14988_/A vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_177_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19225_ _26826_/Q _26794_/Q _26762_/Q _26730_/Q _19203_/X _19111_/X vssd1 vssd1 vccd1
+ vccd1 _19226_/B sky130_fd_sc_hd__mux4_1
X_16437_ _16460_/B vssd1 vssd1 vccd1 vccd1 _16779_/A sky130_fd_sc_hd__clkbuf_2
X_13649_ _13649_/A vssd1 vssd1 vccd1 vccd1 _13661_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_176_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19156_ _26823_/Q _26791_/Q _26759_/Q _26727_/Q _19039_/X _19111_/X vssd1 vssd1 vccd1
+ vccd1 _19157_/B sky130_fd_sc_hd__mux4_1
XFILLER_118_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16368_ _16745_/A vssd1 vssd1 vccd1 vccd1 _16744_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18107_ _26692_/Q _26660_/Q _26628_/Q _26596_/Q _18036_/X _18106_/X vssd1 vssd1 vccd1
+ vccd1 _18108_/A sky130_fd_sc_hd__mux4_1
XFILLER_118_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15319_ _15319_/A vssd1 vssd1 vccd1 vccd1 _15328_/S sky130_fd_sc_hd__clkbuf_2
X_19087_ _19227_/A vssd1 vssd1 vccd1 vccd1 _19087_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16299_ _16296_/X _16297_/Y _16298_/X _16109_/A vssd1 vssd1 vccd1 vccd1 _16648_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18038_ _18038_/A _17978_/X vssd1 vssd1 vccd1 vccd1 _18038_/X sky130_fd_sc_hd__or2b_1
XFILLER_160_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20000_ _19988_/X _19989_/X _19990_/X _19991_/X _19994_/X _19997_/X vssd1 vssd1 vccd1
+ vccd1 _20001_/A sky130_fd_sc_hd__mux4_1
XFILLER_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19989_ _19989_/A vssd1 vssd1 vccd1 vccd1 _19989_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21951_ _21999_/A vssd1 vssd1 vccd1 vccd1 _21951_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _20902_/A vssd1 vssd1 vccd1 vccd1 _20902_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24670_ _27586_/Q _24660_/X _24669_/X _24663_/X vssd1 vssd1 vccd1 vccd1 _27586_/D
+ sky130_fd_sc_hd__o211a_1
X_21882_ _21914_/A vssd1 vssd1 vccd1 vccd1 _21882_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23621_ _23624_/A _23621_/B vssd1 vssd1 vccd1 vccd1 _23622_/A sky130_fd_sc_hd__and2_1
X_20833_ _20865_/A vssd1 vssd1 vccd1 vccd1 _20833_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26340_ _20503_/X _26340_/D vssd1 vssd1 vccd1 vccd1 _26340_/Q sky130_fd_sc_hd__dfxtp_1
X_23552_ _23552_/A vssd1 vssd1 vccd1 vccd1 _27206_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20764_ _20754_/X _20755_/X _20756_/X _20757_/X _20758_/X _20759_/X vssd1 vssd1 vccd1
+ vccd1 _20765_/A sky130_fd_sc_hd__mux4_1
XFILLER_161_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22503_ _22519_/A vssd1 vssd1 vccd1 vccd1 _22503_/X sky130_fd_sc_hd__clkbuf_1
X_26271_ _20259_/X _26271_/D vssd1 vssd1 vccd1 vccd1 _26271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20695_ _20695_/A vssd1 vssd1 vccd1 vccd1 _20695_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23483_ _27186_/Q _23483_/B vssd1 vssd1 vccd1 vccd1 _23483_/X sky130_fd_sc_hd__or2_1
XFILLER_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_28010_ _28010_/A _15969_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
XFILLER_149_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25222_ _27703_/Q _25184_/X _25221_/Y _25214_/X vssd1 vssd1 vccd1 vccd1 _27703_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22434_ _22434_/A vssd1 vssd1 vccd1 vccd1 _22434_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25153_ _27525_/Q _27493_/Q vssd1 vssd1 vccd1 vccd1 _25155_/A sky130_fd_sc_hd__and2_1
X_22365_ _22451_/A vssd1 vssd1 vccd1 vccd1 _22433_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_202_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24104_ _27400_/Q _24106_/B vssd1 vssd1 vccd1 vccd1 _24105_/A sky130_fd_sc_hd__and2_1
X_21316_ _21316_/A vssd1 vssd1 vccd1 vccd1 _21316_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22296_ _22296_/A vssd1 vssd1 vccd1 vccd1 _22296_/X sky130_fd_sc_hd__clkbuf_1
X_25084_ _25084_/A vssd1 vssd1 vccd1 vccd1 _27684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_514 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24035_ _23990_/X _24033_/X _24034_/X _24005_/X vssd1 vssd1 vccd1 vccd1 _27300_/D
+ sky130_fd_sc_hd__o211a_1
X_21247_ _21231_/X _21234_/X _21237_/X _21240_/X _21241_/X _21242_/X vssd1 vssd1 vccd1
+ vccd1 _21248_/A sky130_fd_sc_hd__mux4_1
XFILLER_81_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_453 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_21178_ _21178_/A vssd1 vssd1 vccd1 vccd1 _21178_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20129_ _20129_/A vssd1 vssd1 vccd1 vccd1 _20129_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25986_ _25986_/CLK _25986_/D vssd1 vssd1 vccd1 vccd1 _25986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27725_ _27735_/CLK _27725_/D vssd1 vssd1 vccd1 vccd1 _27725_/Q sky130_fd_sc_hd__dfxtp_1
X_12951_ _12951_/A vssd1 vssd1 vccd1 vccd1 _27820_/D sky130_fd_sc_hd__clkbuf_1
X_24937_ _24937_/A _24937_/B vssd1 vssd1 vccd1 vccd1 _24937_/Y sky130_fd_sc_hd__nand2_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27656_ _27658_/CLK _27656_/D vssd1 vssd1 vccd1 vccd1 _27656_/Q sky130_fd_sc_hd__dfxtp_1
X_15670_ _13172_/X _26149_/Q _15678_/S vssd1 vssd1 vccd1 vccd1 _15671_/A sky130_fd_sc_hd__mux2_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _14497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24868_ _24862_/A _24867_/C _27763_/Q vssd1 vssd1 vccd1 vccd1 _24869_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_211 _14511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _14795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26607_ _21438_/X _26607_/D vssd1 vssd1 vccd1 vccd1 _26607_/Q sky130_fd_sc_hd__dfxtp_1
X_14621_ _26586_/Q _14615_/X _14542_/B _14620_/Y vssd1 vssd1 vccd1 vccd1 _26586_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _17321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23819_ _25918_/Q _25984_/Q _25817_/Q _26016_/Q _23804_/X _23786_/X vssd1 vssd1 vccd1
+ vccd1 _23819_/X sky130_fd_sc_hd__mux4_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _25641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_27587_ _27587_/CLK _27587_/D vssd1 vssd1 vccd1 vccd1 _27587_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _26815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24799_ _24941_/A vssd1 vssd1 vccd1 vccd1 _24800_/A sky130_fd_sc_hd__inv_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_751 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17338_/X _17340_/B vssd1 vssd1 vccd1 vccd1 _17340_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_277 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14552_ _14552_/A vssd1 vssd1 vccd1 vccd1 _14605_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_26538_ _21192_/X _26538_/D vssd1 vssd1 vccd1 vccd1 _26538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_288 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ _13897_/A _13517_/B vssd1 vssd1 vccd1 vccd1 _13503_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17271_ _17238_/X _17265_/X _17268_/X _17270_/X vssd1 vssd1 vccd1 vccd1 _17271_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _15745_/A _14483_/B vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26469_ _20952_/X _26469_/D vssd1 vssd1 vccd1 vccd1 _26469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19010_ _19004_/X _19006_/X _19009_/X _18866_/X _18987_/X vssd1 vssd1 vccd1 vccd1
+ _19011_/C sky130_fd_sc_hd__a221o_1
XFILLER_186_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16222_ _27381_/Q vssd1 vssd1 vccd1 vccd1 _23033_/A sky130_fd_sc_hd__inv_2
XFILLER_201_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13434_ _26969_/Q _13423_/X _13429_/X _13433_/Y vssd1 vssd1 vccd1 vccd1 _26969_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ _27398_/Q _16297_/B vssd1 vssd1 vccd1 vccd1 _16153_/Y sky130_fd_sc_hd__nand2_1
X_13365_ _13365_/A vssd1 vssd1 vccd1 vccd1 _26988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ _14791_/X _26400_/Q _15112_/S vssd1 vssd1 vccd1 vccd1 _15105_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16084_ _16084_/A vssd1 vssd1 vccd1 vccd1 _16699_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_170_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13296_ _27012_/Q _13179_/X _13302_/S vssd1 vssd1 vccd1 vccd1 _13297_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15035_ _26430_/Q _15028_/X _15029_/X _15034_/Y vssd1 vssd1 vccd1 vccd1 _26430_/D
+ sky130_fd_sc_hd__a31o_1
X_19912_ _19898_/X _19899_/X _19900_/X _19901_/X _19903_/X _19905_/X vssd1 vssd1 vccd1
+ vccd1 _19913_/A sky130_fd_sc_hd__mux4_1
XFILLER_5_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19843_ _19843_/A vssd1 vssd1 vccd1 vccd1 _19843_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19774_ _19764_/X _19765_/X _19766_/X _19767_/X _19768_/X _19769_/X vssd1 vssd1 vccd1
+ vccd1 _19775_/A sky130_fd_sc_hd__mux4_1
X_16986_ input35/X vssd1 vssd1 vccd1 vccd1 _17380_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18725_ _18725_/A vssd1 vssd1 vccd1 vccd1 _26024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15937_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15937_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18656_ _18656_/A vssd1 vssd1 vccd1 vccd1 _25993_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15868_ _15868_/A vssd1 vssd1 vccd1 vccd1 _15868_/Y sky130_fd_sc_hd__inv_2
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14819_ _14819_/A vssd1 vssd1 vccd1 vccd1 _26520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17607_ _17607_/A vssd1 vssd1 vccd1 vccd1 _25876_/D sky130_fd_sc_hd__clkbuf_1
X_18587_ _18605_/A vssd1 vssd1 vccd1 vccd1 _25434_/A sky130_fd_sc_hd__buf_2
X_15799_ _13094_/X _26099_/Q _15805_/S vssd1 vssd1 vccd1 vccd1 _15800_/A sky130_fd_sc_hd__mux2_1
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17538_ _17434_/X _25846_/Q _17540_/S vssd1 vssd1 vccd1 vccd1 _17539_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17469_ _27422_/Q vssd1 vssd1 vccd1 vccd1 _17469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19208_ _19208_/A vssd1 vssd1 vccd1 vccd1 _19208_/X sky130_fd_sc_hd__buf_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater80 _27427_/CLK vssd1 vssd1 vccd1 vccd1 _27437_/CLK sky130_fd_sc_hd__clkbuf_1
X_20480_ _20512_/A vssd1 vssd1 vccd1 vccd1 _20480_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater91 _25895_/CLK vssd1 vssd1 vccd1 vccd1 _27849_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_186_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19139_ _19393_/A vssd1 vssd1 vccd1 vccd1 _19139_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22150_ _22150_/A vssd1 vssd1 vccd1 vccd1 _22150_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21101_ _21093_/X _21094_/X _21095_/X _21096_/X _21097_/X _21098_/X vssd1 vssd1 vccd1
+ vccd1 _21102_/A sky130_fd_sc_hd__mux4_1
XFILLER_195_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22081_ _22067_/X _22068_/X _22069_/X _22070_/X _22071_/X _22072_/X vssd1 vssd1 vccd1
+ vccd1 _22082_/A sky130_fd_sc_hd__mux4_1
XFILLER_172_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21032_ _21032_/A vssd1 vssd1 vccd1 vccd1 _21032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25840_ _26039_/CLK _25840_/D vssd1 vssd1 vccd1 vccd1 _25840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25771_ _17472_/X _27841_/Q _25779_/S vssd1 vssd1 vccd1 vccd1 _25772_/A sky130_fd_sc_hd__mux2_1
X_22983_ _22974_/X _22976_/X _22978_/X _22980_/X _22981_/X _22982_/X vssd1 vssd1 vccd1
+ vccd1 _22984_/A sky130_fd_sc_hd__mux4_1
X_27510_ _27511_/CLK _27510_/D vssd1 vssd1 vccd1 vccd1 _27510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24722_ _27605_/Q _24714_/X _24721_/X _24717_/X vssd1 vssd1 vccd1 vccd1 _27605_/D
+ sky130_fd_sc_hd__o211a_1
X_21934_ _21999_/A vssd1 vssd1 vccd1 vccd1 _21934_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27441_ _27442_/CLK _27441_/D vssd1 vssd1 vccd1 vccd1 _27441_/Q sky130_fd_sc_hd__dfxtp_1
X_24653_ _27579_/Q _24643_/X _24652_/X _24650_/X vssd1 vssd1 vccd1 vccd1 _27579_/D
+ sky130_fd_sc_hd__o211a_1
X_21865_ _21913_/A vssd1 vssd1 vccd1 vccd1 _21865_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23604_ _24947_/A _27221_/Q _23616_/S vssd1 vssd1 vccd1 vccd1 _23605_/B sky130_fd_sc_hd__mux2_1
XFILLER_179_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20816_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20816_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27372_ _27372_/CLK _27372_/D vssd1 vssd1 vccd1 vccd1 _27372_/Q sky130_fd_sc_hd__dfxtp_1
X_24584_ _24584_/A vssd1 vssd1 vccd1 vccd1 _27552_/D sky130_fd_sc_hd__clkbuf_1
X_21796_ _21828_/A vssd1 vssd1 vccd1 vccd1 _21796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_169_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26323_ _20441_/X _26323_/D vssd1 vssd1 vccd1 vccd1 _26323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23535_ _23535_/A vssd1 vssd1 vccd1 vccd1 _27201_/D sky130_fd_sc_hd__clkbuf_1
X_20747_ _20747_/A vssd1 vssd1 vccd1 vccd1 _20747_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26254_ _20199_/X _26254_/D vssd1 vssd1 vccd1 vccd1 _26254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23466_ input17/X _23455_/X _23465_/X _23461_/X vssd1 vssd1 vccd1 vccd1 _27179_/D
+ sky130_fd_sc_hd__o211a_1
X_20678_ _20668_/X _20669_/X _20670_/X _20671_/X _20672_/X _20673_/X vssd1 vssd1 vccd1
+ vccd1 _20679_/A sky130_fd_sc_hd__mux4_1
XFILLER_177_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25205_ _25205_/A _25205_/B vssd1 vssd1 vccd1 vccd1 _25206_/B sky130_fd_sc_hd__xnor2_1
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22417_ _22433_/A vssd1 vssd1 vccd1 vccd1 _22417_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_534 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26185_ _19963_/X _26185_/D vssd1 vssd1 vccd1 vccd1 _26185_/Q sky130_fd_sc_hd__dfxtp_1
X_23397_ _27772_/Q vssd1 vssd1 vccd1 vccd1 _24782_/A sky130_fd_sc_hd__inv_2
XFILLER_195_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _16252_/A vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__buf_2
X_25136_ _25136_/A _25149_/A vssd1 vssd1 vccd1 vccd1 _25138_/A sky130_fd_sc_hd__or2b_1
XFILLER_100_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22348_ _22348_/A vssd1 vssd1 vccd1 vccd1 _22348_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_152_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25067_ _27973_/A _25066_/X _25067_/S vssd1 vssd1 vccd1 vccd1 _25068_/A sky130_fd_sc_hd__mux2_1
X_13081_ _13081_/A vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__clkbuf_4
X_22279_ _22451_/A vssd1 vssd1 vccd1 vccd1 _22347_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24018_ _27093_/Q _27125_/Q _24032_/S vssd1 vssd1 vccd1 vccd1 _24018_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _16800_/A _16834_/X _16839_/X vssd1 vssd1 vccd1 vccd1 _16840_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16771_ _16728_/X _16767_/Y _16768_/X _16780_/A _16770_/Y vssd1 vssd1 vccd1 vccd1
+ _16776_/A sky130_fd_sc_hd__a2111o_1
X_13983_ _14038_/A vssd1 vssd1 vccd1 vccd1 _13983_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25969_ _25969_/CLK _25969_/D vssd1 vssd1 vccd1 vccd1 _25969_/Q sky130_fd_sc_hd__dfxtp_1
X_15722_ _15761_/A vssd1 vssd1 vccd1 vccd1 _15732_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_18510_ _18510_/A vssd1 vssd1 vccd1 vccd1 _25971_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27708_ _27709_/CLK _27708_/D vssd1 vssd1 vccd1 vccd1 _27708_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ input2/X _12934_/B vssd1 vssd1 vccd1 vccd1 _12935_/A sky130_fd_sc_hd__and2b_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _26421_/Q _26389_/Q _26357_/Q _26325_/Q _19465_/X _19399_/X vssd1 vssd1 vccd1
+ vccd1 _19490_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _26418_/Q _26386_/Q _26354_/Q _26322_/Q _18305_/X _18329_/X vssd1 vssd1 vccd1
+ vccd1 _18441_/X sky130_fd_sc_hd__mux4_1
X_15653_ _15653_/A vssd1 vssd1 vccd1 vccd1 _26157_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27639_ _27720_/CLK _27639_/D vssd1 vssd1 vccd1 vccd1 _27639_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _26593_/Q _14602_/X _14592_/X _14603_/Y vssd1 vssd1 vccd1 vccd1 _26593_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18489_/A vssd1 vssd1 vccd1 vccd1 _18372_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15584_ _26187_/Q _14756_/A _15584_/S vssd1 vssd1 vccd1 vccd1 _15585_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _27220_/Q _17321_/X _17367_/S vssd1 vssd1 vccd1 vccd1 _17324_/A sky130_fd_sc_hd__mux2_1
X_14535_ _14552_/A vssd1 vssd1 vccd1 vccd1 _14620_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17254_ _25932_/Q _25998_/Q _17254_/S vssd1 vssd1 vccd1 vccd1 _17255_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ _26637_/Q _14460_/X _14455_/X _14465_/Y vssd1 vssd1 vccd1 vccd1 _26637_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16205_ _16205_/A vssd1 vssd1 vccd1 vccd1 _16235_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13417_ _14807_/A vssd1 vssd1 vccd1 vccd1 _13417_/X sky130_fd_sc_hd__buf_4
XFILLER_174_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17185_ _17307_/A vssd1 vssd1 vccd1 vccd1 _17234_/S sky130_fd_sc_hd__clkbuf_2
X_14397_ _26657_/Q _14392_/X _14385_/X _14396_/Y vssd1 vssd1 vccd1 vccd1 _26657_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_155_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ _16136_/A _16240_/C vssd1 vssd1 vccd1 vccd1 _16137_/A sky130_fd_sc_hd__nor2_1
X_13348_ _26993_/Q _13347_/X _13351_/S vssd1 vssd1 vccd1 vccd1 _13349_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16067_ _16313_/B _16313_/C _16457_/B vssd1 vssd1 vccd1 vccd1 _16067_/X sky130_fd_sc_hd__a21o_1
X_13279_ _13279_/A vssd1 vssd1 vccd1 vccd1 _27020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15018_ _26437_/Q _15015_/X _15016_/X _15017_/Y vssd1 vssd1 vccd1 vccd1 _26437_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_570 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19826_ _19812_/X _19813_/X _19814_/X _19815_/X _19817_/X _19819_/X vssd1 vssd1 vccd1
+ vccd1 _19827_/A sky130_fd_sc_hd__mux4_1
XFILLER_151_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19757_ _19757_/A vssd1 vssd1 vccd1 vccd1 _19757_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16969_ _24511_/A vssd1 vssd1 vccd1 vccd1 _24435_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18708_ _18708_/A vssd1 vssd1 vccd1 vccd1 _26016_/D sky130_fd_sc_hd__clkbuf_1
X_19688_ _19678_/X _19679_/X _19680_/X _19681_/X _19682_/X _19683_/X vssd1 vssd1 vccd1
+ vccd1 _19689_/A sky130_fd_sc_hd__mux4_1
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _25986_/Q _17702_/X _18641_/S vssd1 vssd1 vccd1 vccd1 _18640_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21650_ _21650_/A vssd1 vssd1 vccd1 vccd1 _21650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20601_ _20601_/A vssd1 vssd1 vccd1 vccd1 _20601_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21581_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21648_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23320_ _23320_/A _23320_/B _23320_/C _23319_/X vssd1 vssd1 vccd1 vccd1 _23321_/D
+ sky130_fd_sc_hd__or4b_1
X_20532_ _20704_/A vssd1 vssd1 vccd1 vccd1 _20599_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23251_ _23251_/A vssd1 vssd1 vccd1 vccd1 _27160_/D sky130_fd_sc_hd__clkbuf_1
X_20463_ _20463_/A vssd1 vssd1 vccd1 vccd1 _20463_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22202_ _22250_/A vssd1 vssd1 vccd1 vccd1 _22202_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_23182_ _27379_/Q _23182_/B _25735_/C vssd1 vssd1 vccd1 vccd1 _23239_/A sky130_fd_sc_hd__or3_4
X_20394_ _20426_/A vssd1 vssd1 vccd1 vccd1 _20394_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22133_ _22125_/X _22126_/X _22127_/X _22128_/X _22129_/X _22130_/X vssd1 vssd1 vccd1
+ vccd1 _22134_/A sky130_fd_sc_hd__mux4_1
XFILLER_160_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27990_ _27990_/A _15892_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
X_26941_ _22602_/X _26941_/D vssd1 vssd1 vccd1 vccd1 _26941_/Q sky130_fd_sc_hd__dfxtp_1
X_22064_ _22064_/A vssd1 vssd1 vccd1 vccd1 _22064_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21015_ _21007_/X _21008_/X _21009_/X _21010_/X _21011_/X _21012_/X vssd1 vssd1 vccd1
+ vccd1 _21016_/A sky130_fd_sc_hd__mux4_1
X_26872_ _22360_/X _26872_/D vssd1 vssd1 vccd1 vccd1 _26872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25823_ _26022_/CLK _25823_/D vssd1 vssd1 vccd1 vccd1 _25823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25754_ _25754_/A vssd1 vssd1 vccd1 vccd1 _27833_/D sky130_fd_sc_hd__clkbuf_1
X_22966_ _22966_/A vssd1 vssd1 vccd1 vccd1 _22966_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24705_ _27183_/Q _24711_/B vssd1 vssd1 vccd1 vccd1 _24705_/X sky130_fd_sc_hd__or2_1
X_21917_ _22089_/A vssd1 vssd1 vccd1 vccd1 _21986_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25685_ _25673_/X _25674_/X _25675_/X _25676_/X _25677_/X _25678_/X vssd1 vssd1 vccd1
+ vccd1 _25686_/A sky130_fd_sc_hd__mux4_1
X_22897_ _22888_/X _22890_/X _22892_/X _22894_/X _22895_/X _22896_/X vssd1 vssd1 vccd1
+ vccd1 _22898_/A sky130_fd_sc_hd__mux4_1
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27424_ _27425_/CLK _27424_/D vssd1 vssd1 vccd1 vccd1 _27424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24636_ _24636_/A _24636_/B _24636_/C vssd1 vssd1 vccd1 vccd1 _24637_/A sky130_fd_sc_hd__and3_1
XFILLER_71_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21848_ _21913_/A vssd1 vssd1 vccd1 vccd1 _21848_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27355_ _27365_/CLK _27355_/D vssd1 vssd1 vccd1 vccd1 _27355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24567_ _24589_/A vssd1 vssd1 vccd1 vccd1 _24576_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_21779_ _21827_/A vssd1 vssd1 vccd1 vccd1 _21779_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14320_ _14408_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14320_/Y sky130_fd_sc_hd__nor2_1
X_26306_ _20385_/X _26306_/D vssd1 vssd1 vccd1 vccd1 _26306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23518_ _23526_/A _23518_/B vssd1 vssd1 vccd1 vccd1 _23519_/A sky130_fd_sc_hd__and2_1
XFILLER_196_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27286_ _27288_/CLK _27286_/D vssd1 vssd1 vccd1 vccd1 _27286_/Q sky130_fd_sc_hd__dfxtp_1
X_24498_ _27586_/Q _24505_/B vssd1 vssd1 vccd1 vccd1 _24498_/X sky130_fd_sc_hd__or2_1
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14251_ _14304_/A vssd1 vssd1 vccd1 vccd1 _14263_/B sky130_fd_sc_hd__clkbuf_2
X_26237_ _20141_/X _26237_/D vssd1 vssd1 vccd1 vccd1 _26237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_459 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23449_ _27173_/Q _23456_/B vssd1 vssd1 vccd1 vccd1 _23449_/X sky130_fd_sc_hd__or2_1
X_13202_ _27341_/Q _13017_/A _13025_/A _27309_/Q _13201_/X vssd1 vssd1 vccd1 vccd1
+ _16212_/A sky130_fd_sc_hd__a221o_1
X_14182_ _14359_/A _14187_/B vssd1 vssd1 vccd1 vccd1 _14182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26168_ _19895_/X _26168_/D vssd1 vssd1 vccd1 vccd1 _26168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25119_ _27521_/Q _27489_/Q vssd1 vssd1 vccd1 vccd1 _25119_/X sky130_fd_sc_hd__and2_1
X_13133_ _14753_/A vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__buf_2
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26099_ _19657_/X _26099_/D vssd1 vssd1 vccd1 vccd1 _26099_/Q sky130_fd_sc_hd__dfxtp_1
X_18990_ _18990_/A vssd1 vssd1 vccd1 vccd1 _26047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_180_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_653 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _17830_/X _17938_/X _17940_/X vssd1 vssd1 vccd1 vccd1 _17941_/X sky130_fd_sc_hd__o21a_1
X_13064_ _13102_/A vssd1 vssd1 vccd1 vccd1 _13064_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_133_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17872_ _17872_/A _17827_/X vssd1 vssd1 vccd1 vccd1 _17872_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater209 _27417_/CLK vssd1 vssd1 vccd1 vccd1 _26018_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19611_ _19605_/X _19606_/X _19607_/X _19608_/X _19609_/X _19610_/X vssd1 vssd1 vccd1
+ vccd1 _19612_/A sky130_fd_sc_hd__mux4_1
X_16823_ _16534_/A _16535_/A _16804_/Y _16822_/X vssd1 vssd1 vccd1 vccd1 _16823_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19542_ _19560_/A _19542_/B vssd1 vssd1 vccd1 vccd1 _19542_/X sky130_fd_sc_hd__or2_1
X_13966_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14346_/A sky130_fd_sc_hd__buf_2
X_16754_ _16754_/A vssd1 vssd1 vccd1 vccd1 _16754_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15705_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19473_ _19473_/A vssd1 vssd1 vccd1 vccd1 _19567_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16685_ _16450_/A _16450_/B _16684_/X vssd1 vssd1 vccd1 vccd1 _16686_/B sky130_fd_sc_hd__a21oi_1
X_13897_ _13897_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _18424_/A vssd1 vssd1 vccd1 vccd1 _25967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15636_ _15693_/S vssd1 vssd1 vccd1 vccd1 _15645_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18355_ _27814_/Q _26575_/Q _26447_/Q _26127_/Q _18242_/X _18267_/X vssd1 vssd1 vccd1
+ vccd1 _18355_/X sky130_fd_sc_hd__mux4_2
X_15567_ _26195_/Q _14731_/A _15573_/S vssd1 vssd1 vccd1 vccd1 _15568_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17306_ _17299_/X _17300_/X _17302_/X _17305_/X vssd1 vssd1 vccd1 vccd1 _17306_/X
+ sky130_fd_sc_hd__o22a_1
X_14518_ _14518_/A vssd1 vssd1 vccd1 vccd1 _15771_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18286_ _18278_/X _18281_/X _18284_/X _18285_/X _18238_/X vssd1 vssd1 vccd1 vccd1
+ _18287_/C sky130_fd_sc_hd__a221o_1
X_15498_ _15498_/A vssd1 vssd1 vccd1 vccd1 _26226_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_175_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14465_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_17237_ _17237_/A vssd1 vssd1 vccd1 vccd1 _27934_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_163_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _17155_/X _17168_/B vssd1 vssd1 vccd1 vccd1 _17168_/X sky130_fd_sc_hd__and2b_1
XFILLER_7_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16119_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16119_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17099_ _17057_/X _17097_/X _17098_/X vssd1 vssd1 vccd1 vccd1 _17099_/X sky130_fd_sc_hd__a21bo_1
XFILLER_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_432 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19809_ _19809_/A vssd1 vssd1 vccd1 vccd1 _19809_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22820_ _22820_/A vssd1 vssd1 vccd1 vccd1 _22820_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22751_ _22783_/A vssd1 vssd1 vccd1 vccd1 _22751_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21702_ _21702_/A vssd1 vssd1 vccd1 vccd1 _21702_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25470_ _25560_/A vssd1 vssd1 vccd1 vccd1 _25470_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_198_849 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22682_ _22698_/A vssd1 vssd1 vccd1 vccd1 _22682_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_201_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24421_ _24421_/A vssd1 vssd1 vccd1 vccd1 _27489_/D sky130_fd_sc_hd__clkbuf_1
X_21633_ _21649_/A vssd1 vssd1 vccd1 vccd1 _21633_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27140_ _27140_/CLK _27140_/D vssd1 vssd1 vccd1 vccd1 _27140_/Q sky130_fd_sc_hd__dfxtp_1
X_24352_ _24363_/A vssd1 vssd1 vccd1 vccd1 _24361_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_178_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21564_ _21564_/A vssd1 vssd1 vccd1 vccd1 _21564_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23303_ _27735_/Q _23296_/Y _23302_/Y input64/X vssd1 vssd1 vccd1 vccd1 _23303_/Y
+ sky130_fd_sc_hd__o22ai_1
X_20515_ _20515_/A vssd1 vssd1 vccd1 vccd1 _20515_/X sky130_fd_sc_hd__clkbuf_1
X_27071_ _27103_/CLK _27071_/D vssd1 vssd1 vccd1 vccd1 _27071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24283_ _16162_/Y _16445_/X _24269_/X vssd1 vssd1 vccd1 vccd1 _27419_/D sky130_fd_sc_hd__o21a_1
XFILLER_165_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21495_ _21581_/A vssd1 vssd1 vccd1 vccd1 _21562_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26022_ _26022_/CLK _26022_/D vssd1 vssd1 vccd1 vccd1 _26022_/Q sky130_fd_sc_hd__dfxtp_1
X_23234_ _23234_/A vssd1 vssd1 vccd1 vccd1 _27152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20446_ _20704_/A vssd1 vssd1 vccd1 vccd1 _20513_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23165_ _27122_/Q _17753_/X _23165_/S vssd1 vssd1 vccd1 vccd1 _23166_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20377_ _20425_/A vssd1 vssd1 vccd1 vccd1 _20377_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22116_ _22116_/A vssd1 vssd1 vccd1 vccd1 _22116_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_23096_ _23096_/A vssd1 vssd1 vccd1 vccd1 _27091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27973_ _27973_/A _15937_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_645 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22047_ _22035_/X _22036_/X _22037_/X _22038_/X _22039_/X _22040_/X vssd1 vssd1 vccd1
+ vccd1 _22048_/A sky130_fd_sc_hd__mux4_1
X_26924_ _22536_/X _26924_/D vssd1 vssd1 vccd1 vccd1 _26924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26855_ _22306_/X _26855_/D vssd1 vssd1 vccd1 vccd1 _26855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_424 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _13833_/A vssd1 vssd1 vccd1 vccd1 _13820_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25806_ _25806_/A vssd1 vssd1 vccd1 vccd1 _27857_/D sky130_fd_sc_hd__clkbuf_1
X_26786_ _22060_/X _26786_/D vssd1 vssd1 vccd1 vccd1 _26786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23998_ _27091_/Q _27123_/Q _24032_/S vssd1 vssd1 vccd1 vccd1 _23998_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _13930_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13751_/Y sky130_fd_sc_hd__nor2_1
X_25737_ _25805_/S vssd1 vssd1 vccd1 vccd1 _25746_/S sky130_fd_sc_hd__clkbuf_2
X_22949_ _22939_/X _22940_/X _22941_/X _22942_/X _22943_/X _22944_/X vssd1 vssd1 vccd1
+ vccd1 _22950_/A sky130_fd_sc_hd__mux4_1
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_816 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16470_ _16470_/A vssd1 vssd1 vccd1 vccd1 _16778_/B sky130_fd_sc_hd__inv_2
X_13682_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13682_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25668_ _25668_/A vssd1 vssd1 vccd1 vccd1 _25668_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15421_ _26260_/Q _13337_/X _15429_/S vssd1 vssd1 vccd1 vccd1 _15422_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24619_ _24619_/A vssd1 vssd1 vccd1 vccd1 _27568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27407_ _27407_/CLK _27407_/D vssd1 vssd1 vccd1 vccd1 _27407_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25599_ _25438_/X _25336_/B _25598_/X _18591_/X vssd1 vssd1 vccd1 vccd1 _25599_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_1163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15352_ _15352_/A vssd1 vssd1 vccd1 vccd1 _26291_/D sky130_fd_sc_hd__clkbuf_1
X_18140_ _18020_/X _18139_/X _18070_/X vssd1 vssd1 vccd1 vccd1 _18140_/X sky130_fd_sc_hd__o21a_1
X_27338_ _27338_/CLK _27338_/D vssd1 vssd1 vccd1 vccd1 _27338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14303_ _26691_/Q _14296_/X _14297_/X _14302_/Y vssd1 vssd1 vccd1 vccd1 _26691_/D
+ sky130_fd_sc_hd__a31o_1
X_18071_ _18020_/X _18069_/X _18070_/X vssd1 vssd1 vccd1 vccd1 _18071_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15283_ _15283_/A vssd1 vssd1 vccd1 vccd1 _26321_/D sky130_fd_sc_hd__clkbuf_1
X_27269_ _27335_/CLK _27269_/D vssd1 vssd1 vccd1 vccd1 _27269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17022_ _16998_/X _17021_/X _17299_/A vssd1 vssd1 vccd1 vccd1 _17022_/X sky130_fd_sc_hd__a21bo_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14234_ _14412_/A _14234_/B vssd1 vssd1 vccd1 vccd1 _14234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14165_ _26741_/Q _14157_/X _14151_/X _14164_/Y vssd1 vssd1 vccd1 vccd1 _26741_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _14743_/A vssd1 vssd1 vccd1 vccd1 _13116_/X sky130_fd_sc_hd__buf_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14361_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14096_/Y sky130_fd_sc_hd__nor2_1
X_18973_ _26943_/Q _26911_/Q _26879_/Q _26847_/Q _18875_/X _18972_/X vssd1 vssd1 vccd1
+ vccd1 _18973_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13425_/A _13672_/A _27265_/Q _13244_/B vssd1 vssd1 vccd1 vccd1 _15551_/A
+ sky130_fd_sc_hd__nand4_4
X_17924_ _17924_/A vssd1 vssd1 vccd1 vccd1 _18437_/A sky130_fd_sc_hd__buf_2
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17855_ _18489_/A vssd1 vssd1 vccd1 vccd1 _18238_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _16801_/X _16802_/Y _16803_/Y _16804_/Y _16805_/Y vssd1 vssd1 vccd1 vccd1
+ _16806_/X sky130_fd_sc_hd__a2111o_1
XFILLER_54_608 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17786_ _27793_/Q _26554_/Q _26426_/Q _26106_/Q _17782_/X _17785_/X vssd1 vssd1 vccd1
+ vccd1 _17786_/X sky130_fd_sc_hd__mux4_2
X_14998_ _26444_/Q _14988_/X _14989_/X _14997_/Y vssd1 vssd1 vccd1 vccd1 _26444_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19525_ _26295_/Q _26263_/Q _26231_/Q _26199_/Q _19441_/X _19486_/X vssd1 vssd1 vccd1
+ vccd1 _19525_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16737_ _16737_/A _16737_/B _16737_/C vssd1 vssd1 vccd1 vccd1 _16737_/X sky130_fd_sc_hd__and3_1
X_13949_ _14005_/A vssd1 vssd1 vccd1 vccd1 _13949_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_449 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19456_ _26964_/Q _26932_/Q _26900_/Q _26868_/Q _19343_/X _19412_/X vssd1 vssd1 vccd1
+ vccd1 _19456_/X sky130_fd_sc_hd__mux4_1
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668_ _16093_/X _16664_/X _16667_/X _16626_/X vssd1 vssd1 vccd1 vccd1 _24245_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18407_ _26833_/Q _26801_/Q _26769_/Q _26737_/Q _18358_/X _18380_/X vssd1 vssd1 vccd1
+ vccd1 _18407_/X sky130_fd_sc_hd__mux4_2
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _26171_/Q _14807_/A _15621_/S vssd1 vssd1 vccd1 vccd1 _15620_/A sky130_fd_sc_hd__mux2_1
X_19387_ _19387_/A vssd1 vssd1 vccd1 vccd1 _19387_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16599_ _16599_/A _16599_/B vssd1 vssd1 vccd1 vccd1 _16599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18338_ _18020_/A _18337_/X _18014_/A vssd1 vssd1 vccd1 vccd1 _18338_/X sky130_fd_sc_hd__o21a_1
XFILLER_148_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18269_ _18427_/A vssd1 vssd1 vccd1 vccd1 _18269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20300_ _20286_/X _20287_/X _20288_/X _20289_/X _20290_/X _20291_/X vssd1 vssd1 vccd1
+ vccd1 _20301_/A sky130_fd_sc_hd__mux4_1
XFILLER_162_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21280_ _21280_/A vssd1 vssd1 vccd1 vccd1 _21280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20231_ _20231_/A vssd1 vssd1 vccd1 vccd1 _20231_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20162_ _20162_/A vssd1 vssd1 vccd1 vccd1 _20162_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24970_ _24970_/A _24970_/B vssd1 vssd1 vccd1 vccd1 _24970_/Y sky130_fd_sc_hd__nand2_1
X_20093_ _20093_/A vssd1 vssd1 vccd1 vccd1 _20093_/X sky130_fd_sc_hd__clkbuf_1
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23921_ _27843_/Q _27147_/Q _25892_/Q _25860_/Q _23920_/X _23897_/X vssd1 vssd1 vccd1
+ vccd1 _23921_/X sky130_fd_sc_hd__mux4_1
XFILLER_97_582 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26640_ _21552_/X _26640_/D vssd1 vssd1 vccd1 vccd1 _26640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23852_ _23946_/A vssd1 vssd1 vccd1 vccd1 _23852_/X sky130_fd_sc_hd__buf_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_22803_ _22889_/A vssd1 vssd1 vccd1 vccd1 _22870_/A sky130_fd_sc_hd__clkbuf_2
X_26571_ _21314_/X _26571_/D vssd1 vssd1 vccd1 vccd1 _26571_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_438 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23783_ _27068_/Q _23761_/X _23763_/X _27100_/Q _23765_/X vssd1 vssd1 vccd1 vccd1
+ _23783_/X sky130_fd_sc_hd__a221o_1
X_20995_ _21027_/A vssd1 vssd1 vccd1 vccd1 _20995_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25522_ _25552_/A vssd1 vssd1 vccd1 vccd1 _25522_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22734_ _22734_/A vssd1 vssd1 vccd1 vccd1 _22734_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25453_ _25438_/X _25131_/B _25451_/X _25452_/X vssd1 vssd1 vccd1 vccd1 _25453_/X
+ sky130_fd_sc_hd__a211o_1
X_22665_ _22697_/A vssd1 vssd1 vccd1 vccd1 _22665_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_24404_ _24404_/A vssd1 vssd1 vccd1 vccd1 _27481_/D sky130_fd_sc_hd__clkbuf_1
X_21616_ _21648_/A vssd1 vssd1 vccd1 vccd1 _21616_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25384_ _25384_/A vssd1 vssd1 vccd1 vccd1 _27731_/D sky130_fd_sc_hd__clkbuf_1
X_22596_ _22612_/A vssd1 vssd1 vccd1 vccd1 _22596_/X sky130_fd_sc_hd__clkbuf_1
X_27123_ _27123_/CLK _27123_/D vssd1 vssd1 vccd1 vccd1 _27123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24335_ _27551_/Q _24339_/B vssd1 vssd1 vccd1 vccd1 _24336_/A sky130_fd_sc_hd__and2_1
X_21547_ _21563_/A vssd1 vssd1 vccd1 vccd1 _21547_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_407 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27054_ _22992_/X _27054_/D vssd1 vssd1 vccd1 vccd1 _27054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24266_ _25517_/A vssd1 vssd1 vccd1 vccd1 _24267_/A sky130_fd_sc_hd__clkbuf_2
X_21478_ _21478_/A vssd1 vssd1 vccd1 vccd1 _21478_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1041 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26005_ _27149_/CLK _26005_/D vssd1 vssd1 vccd1 vccd1 _26005_/Q sky130_fd_sc_hd__dfxtp_1
X_23217_ _23239_/A vssd1 vssd1 vccd1 vccd1 _23226_/S sky130_fd_sc_hd__clkbuf_2
X_20429_ _20774_/A vssd1 vssd1 vccd1 vccd1 _20500_/A sky130_fd_sc_hd__clkbuf_2
X_24197_ _27754_/Q _25358_/A vssd1 vssd1 vccd1 vccd1 _24238_/A sky130_fd_sc_hd__nor2_1
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23148_ _27114_/Q _17728_/X _23154_/S vssd1 vssd1 vccd1 vccd1 _23149_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_921 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23079_ _27084_/Q _17734_/X _23081_/S vssd1 vssd1 vccd1 vccd1 _23080_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15970_ _15973_/A vssd1 vssd1 vccd1 vccd1 _15970_/Y sky130_fd_sc_hd__inv_2
X_27956_ _27956_/A _15916_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
XFILLER_96_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26907_ _22482_/X _26907_/D vssd1 vssd1 vccd1 vccd1 _26907_/Q sky130_fd_sc_hd__dfxtp_1
X_14921_ _14759_/X _26474_/Q _14929_/S vssd1 vssd1 vccd1 vccd1 _14922_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17640_ _17640_/A vssd1 vssd1 vccd1 vccd1 _25891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26838_ _22242_/X _26838_/D vssd1 vssd1 vccd1 vccd1 _26838_/Q sky130_fd_sc_hd__dfxtp_1
X_14852_ _14852_/A vssd1 vssd1 vccd1 vccd1 _26505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _26860_/Q _13793_/X _13794_/X _13802_/Y vssd1 vssd1 vccd1 vccd1 _26860_/D
+ sky130_fd_sc_hd__a31o_1
X_17571_ _17482_/X _25861_/Q _17573_/S vssd1 vssd1 vccd1 vccd1 _17572_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14783_ _14782_/X _26531_/Q _14789_/S vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26769_ _21996_/X _26769_/D vssd1 vssd1 vccd1 vccd1 _26769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _19304_/X _19306_/X _19309_/X _18895_/A vssd1 vssd1 vccd1 vccd1 _19310_/X
+ sky130_fd_sc_hd__a22o_1
X_13734_ _26885_/Q _13724_/X _13732_/X _13733_/Y vssd1 vssd1 vccd1 vccd1 _26885_/D
+ sky130_fd_sc_hd__a31o_1
X_16522_ _25967_/Q _16412_/X _16521_/X vssd1 vssd1 vccd1 vccd1 _16826_/A sky130_fd_sc_hd__a21oi_4
XFILLER_45_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_460 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19241_ _26410_/Q _26378_/Q _26346_/Q _26314_/Q _19170_/X _19240_/X vssd1 vssd1 vccd1
+ vccd1 _19241_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13665_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16453_ _16453_/A vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A vssd1 vssd1 vccd1 vccd1 _26267_/D sky130_fd_sc_hd__clkbuf_1
X_19172_ _26535_/Q _26503_/Q _26471_/Q _27047_/Q _19102_/X _19148_/X vssd1 vssd1 vccd1
+ vccd1 _19172_/X sky130_fd_sc_hd__mux4_1
X_16384_ _16384_/A vssd1 vssd1 vccd1 vccd1 _16384_/X sky130_fd_sc_hd__clkbuf_2
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13649_/A vssd1 vssd1 vccd1 vccd1 _13608_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15335_ _15335_/A _15551_/B vssd1 vssd1 vccd1 vccd1 _15392_/A sky130_fd_sc_hd__or2_2
X_18123_ _18114_/X _18116_/X _18121_/X _18026_/X _18122_/X vssd1 vssd1 vccd1 vccd1
+ _18124_/C sky130_fd_sc_hd__a221o_1
XFILLER_77_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18054_ _27801_/Q _26562_/Q _26434_/Q _26114_/Q _17920_/X _17949_/X vssd1 vssd1 vccd1
+ vccd1 _18054_/X sky130_fd_sc_hd__mux4_2
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15266_ _15266_/A vssd1 vssd1 vccd1 vccd1 _26329_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_3 _20701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ _26722_/Q _14212_/X _14207_/X _14216_/Y vssd1 vssd1 vccd1 vccd1 _26722_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17005_ _27066_/Q _27098_/Q _17047_/S vssd1 vssd1 vccd1 vccd1 _17005_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15197_ _14718_/X _26359_/Q _15201_/S vssd1 vssd1 vccd1 vccd1 _15198_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14148_ _26746_/Q _14142_/X _14070_/B _14147_/Y vssd1 vssd1 vccd1 vccd1 _26746_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14079_ _14079_/A vssd1 vssd1 vccd1 vccd1 _14133_/A sky130_fd_sc_hd__clkbuf_2
X_18956_ _26270_/Q _26238_/Q _26206_/Q _26174_/Q _18859_/X _18955_/X vssd1 vssd1 vccd1
+ vccd1 _18956_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17907_ _17902_/X _17905_/X _18522_/S vssd1 vssd1 vccd1 vccd1 _17907_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18887_ _19343_/A vssd1 vssd1 vccd1 vccd1 _18887_/X sky130_fd_sc_hd__buf_2
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17838_ _18014_/A vssd1 vssd1 vccd1 vccd1 _17838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17769_ _27437_/Q vssd1 vssd1 vccd1 vccd1 _17769_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19508_ _19485_/X _19507_/X _19488_/X vssd1 vssd1 vccd1 vccd1 _19508_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20780_ _20770_/X _20771_/X _20772_/X _20773_/X _20775_/X _20777_/X vssd1 vssd1 vccd1
+ vccd1 _20781_/A sky130_fd_sc_hd__mux4_1
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _26163_/Q _26099_/Q _27027_/Q _26995_/Q _19326_/X _19348_/X vssd1 vssd1 vccd1
+ vccd1 _19440_/B sky130_fd_sc_hd__mux4_1
XFILLER_23_858 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22450_ _22450_/A vssd1 vssd1 vccd1 vccd1 _22450_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21401_ _21389_/X _21390_/X _21391_/X _21392_/X _21394_/X _21396_/X vssd1 vssd1 vccd1
+ vccd1 _21402_/A sky130_fd_sc_hd__mux4_1
XFILLER_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22381_ _22366_/X _22368_/X _22370_/X _22372_/X _22373_/X _22374_/X vssd1 vssd1 vccd1
+ vccd1 _22382_/A sky130_fd_sc_hd__mux4_1
XFILLER_136_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24120_ _27407_/Q _24128_/B vssd1 vssd1 vccd1 vccd1 _24121_/A sky130_fd_sc_hd__and2_1
XFILLER_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21332_ _21332_/A vssd1 vssd1 vccd1 vccd1 _21332_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24051_ _24051_/A vssd1 vssd1 vccd1 vccd1 _27303_/D sky130_fd_sc_hd__clkbuf_1
X_21263_ _21253_/X _21254_/X _21255_/X _21256_/X _21257_/X _21258_/X vssd1 vssd1 vccd1
+ vccd1 _21264_/A sky130_fd_sc_hd__mux4_1
XFILLER_117_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23002_ _23002_/A vssd1 vssd1 vccd1 vccd1 _23002_/X sky130_fd_sc_hd__clkbuf_1
X_20214_ _20200_/X _20201_/X _20202_/X _20203_/X _20204_/X _20205_/X vssd1 vssd1 vccd1
+ vccd1 _20215_/A sky130_fd_sc_hd__mux4_1
XFILLER_131_410 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21194_ _21194_/A vssd1 vssd1 vccd1 vccd1 _21194_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27810_ _25686_/X _27810_/D vssd1 vssd1 vccd1 vccd1 _27810_/Q sky130_fd_sc_hd__dfxtp_1
X_27951__437 vssd1 vssd1 vccd1 vccd1 _27951__437/HI _27951_/A sky130_fd_sc_hd__conb_1
X_20145_ _20145_/A vssd1 vssd1 vccd1 vccd1 _20145_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_27741_ _27745_/CLK _27741_/D vssd1 vssd1 vccd1 vccd1 _27741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24953_ _27667_/Q _24935_/X _24952_/Y _24938_/X vssd1 vssd1 vccd1 vccd1 _27667_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _20076_/A vssd1 vssd1 vccd1 vccd1 _20076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23904_ _27081_/Q _27113_/Q _23939_/S vssd1 vssd1 vccd1 vccd1 _23904_/X sky130_fd_sc_hd__mux2_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27672_ _27672_/CLK _27672_/D vssd1 vssd1 vccd1 vccd1 _27963_/A sky130_fd_sc_hd__dfxtp_1
X_24884_ _27653_/Q _24861_/X _24883_/Y _24864_/X vssd1 vssd1 vccd1 vccd1 _27653_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater370 _27224_/CLK vssd1 vssd1 vccd1 vccd1 _27677_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater381 _27462_/CLK vssd1 vssd1 vccd1 vccd1 _27563_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26623_ _21490_/X _26623_/D vssd1 vssd1 vccd1 vccd1 _26623_/Q sky130_fd_sc_hd__dfxtp_1
X_23835_ _23929_/A vssd1 vssd1 vccd1 vccd1 _23835_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater392 _27342_/CLK vssd1 vssd1 vccd1 vccd1 _27447_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26554_ _21252_/X _26554_/D vssd1 vssd1 vccd1 vccd1 _26554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23766_ _27066_/Q _23761_/X _23763_/X _27098_/Q _23765_/X vssd1 vssd1 vccd1 vccd1
+ _23766_/X sky130_fd_sc_hd__a221o_1
X_20978_ _21042_/A vssd1 vssd1 vccd1 vccd1 _20978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25505_ _27701_/Q _25479_/X _25480_/X vssd1 vssd1 vccd1 vccd1 _25505_/Y sky130_fd_sc_hd__a21oi_1
X_22717_ _22889_/A vssd1 vssd1 vccd1 vccd1 _22784_/A sky130_fd_sc_hd__buf_2
XFILLER_199_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26485_ _21014_/X _26485_/D vssd1 vssd1 vccd1 vccd1 _26485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_937 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23697_ _27773_/Q _27253_/Q _23705_/S vssd1 vssd1 vccd1 vccd1 _23698_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_25436_ _27691_/Q _25433_/X _25435_/X vssd1 vssd1 vccd1 vccd1 _25436_/Y sky130_fd_sc_hd__a21oi_1
X_13450_ _13529_/A vssd1 vssd1 vccd1 vccd1 _13450_/X sky130_fd_sc_hd__buf_4
X_22648_ _22648_/A vssd1 vssd1 vccd1 vccd1 _22648_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25367_ _27724_/Q input66/X _25369_/S vssd1 vssd1 vccd1 vccd1 _25368_/A sky130_fd_sc_hd__mux2_1
X_13381_ _13381_/A vssd1 vssd1 vccd1 vccd1 _26983_/D sky130_fd_sc_hd__clkbuf_1
X_22579_ _22611_/A vssd1 vssd1 vccd1 vccd1 _22579_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15120_ _15188_/S vssd1 vssd1 vccd1 vccd1 _15129_/S sky130_fd_sc_hd__buf_2
X_24318_ _24318_/A vssd1 vssd1 vccd1 vccd1 _27443_/D sky130_fd_sc_hd__clkbuf_1
X_27106_ _27832_/CLK _27106_/D vssd1 vssd1 vccd1 vccd1 _27106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25298_ _27712_/Q _25263_/X _25296_/Y _25297_/X vssd1 vssd1 vccd1 vccd1 _27712_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27037_ _22934_/X _27037_/D vssd1 vssd1 vccd1 vccd1 _27037_/Q sky130_fd_sc_hd__dfxtp_1
X_15051_ _14715_/X _26424_/Q _15057_/S vssd1 vssd1 vccd1 vccd1 _15052_/A sky130_fd_sc_hd__mux2_1
X_24249_ _24249_/A _24256_/B vssd1 vssd1 vccd1 vccd1 _27396_/D sky130_fd_sc_hd__nor2_1
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ _16495_/A vssd1 vssd1 vccd1 vccd1 _14372_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_421 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18810_ _18926_/A vssd1 vssd1 vccd1 vccd1 _18810_/X sky130_fd_sc_hd__buf_2
XFILLER_96_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19790_ _19780_/X _19781_/X _19782_/X _19783_/X _19784_/X _19785_/X vssd1 vssd1 vccd1
+ vccd1 _19791_/A sky130_fd_sc_hd__mux4_1
X_18741_ _18741_/A vssd1 vssd1 vccd1 vccd1 _26031_/D sky130_fd_sc_hd__clkbuf_1
X_15953_ _15955_/A vssd1 vssd1 vccd1 vccd1 _15953_/Y sky130_fd_sc_hd__inv_2
X_27939_ _27939_/A _15943_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14904_ _14904_/A vssd1 vssd1 vccd1 vccd1 _26482_/D sky130_fd_sc_hd__clkbuf_1
X_18672_ _26001_/Q _17750_/X _18674_/S vssd1 vssd1 vccd1 vccd1 _18673_/A sky130_fd_sc_hd__mux2_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _15887_/A vssd1 vssd1 vccd1 vccd1 _15884_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _17453_/X _25884_/Q _17623_/S vssd1 vssd1 vccd1 vccd1 _17624_/A sky130_fd_sc_hd__mux2_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _26512_/Q _13350_/X _14835_/S vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__mux2_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _17456_/X _25853_/Q _17562_/S vssd1 vssd1 vccd1 vccd1 _17555_/A sky130_fd_sc_hd__mux2_1
XFILLER_189_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14766_ _14766_/A vssd1 vssd1 vccd1 vccd1 _14766_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _16292_/B _16281_/B _16106_/A vssd1 vssd1 vccd1 vccd1 _16506_/B sky130_fd_sc_hd__o21a_1
X_13717_ _26891_/Q _13710_/X _13705_/X _13716_/Y vssd1 vssd1 vccd1 vccd1 _26891_/D
+ sky130_fd_sc_hd__a31o_1
X_17485_ _27427_/Q vssd1 vssd1 vccd1 vccd1 _17485_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _26559_/Q _14685_/X _14693_/X _14696_/Y vssd1 vssd1 vccd1 vccd1 _26559_/D
+ sky130_fd_sc_hd__a31o_1
X_19224_ _19473_/A vssd1 vssd1 vccd1 vccd1 _19362_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16436_ _16769_/B vssd1 vssd1 vccd1 vccd1 _16779_/B sky130_fd_sc_hd__clkbuf_2
X_13648_ _26915_/Q _13639_/X _13642_/X _13647_/Y vssd1 vssd1 vccd1 vccd1 _26915_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19428_/A vssd1 vssd1 vccd1 vccd1 _19250_/A sky130_fd_sc_hd__clkbuf_1
X_13579_ _13792_/A vssd1 vssd1 vccd1 vccd1 _13639_/A sky130_fd_sc_hd__clkbuf_2
X_16367_ _16745_/B vssd1 vssd1 vccd1 vccd1 _16372_/A sky130_fd_sc_hd__inv_2
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18106_ _18408_/A vssd1 vssd1 vccd1 vccd1 _18106_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_191_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15318_ _15318_/A vssd1 vssd1 vccd1 vccd1 _26305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_184_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19086_ _19113_/A _19086_/B vssd1 vssd1 vccd1 vccd1 _19086_/X sky130_fd_sc_hd__or2_1
X_16298_ _16298_/A _16298_/B _16298_/C vssd1 vssd1 vccd1 vccd1 _16298_/X sky130_fd_sc_hd__or3_1
XFILLER_184_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18037_ _26689_/Q _26657_/Q _26625_/Q _26593_/Q _18036_/X _17928_/X vssd1 vssd1 vccd1
+ vccd1 _18038_/A sky130_fd_sc_hd__mux4_2
X_15249_ _15249_/A vssd1 vssd1 vccd1 vccd1 _26336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19988_ _19988_/A vssd1 vssd1 vccd1 vccd1 _19988_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18939_ _19227_/A vssd1 vssd1 vccd1 vccd1 _18939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_1108 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21950_ _21998_/A vssd1 vssd1 vccd1 vccd1 _21950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20901_ _20886_/X _20888_/X _20890_/X _20892_/X _20893_/X _20894_/X vssd1 vssd1 vccd1
+ vccd1 _20902_/A sky130_fd_sc_hd__mux4_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21881_ _21913_/A vssd1 vssd1 vccd1 vccd1 _21881_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23620_ _24965_/A _27225_/Q _23623_/S vssd1 vssd1 vccd1 vccd1 _23621_/B sky130_fd_sc_hd__mux2_1
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20832_ _20864_/A vssd1 vssd1 vccd1 vccd1 _20832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23551_ _23560_/A _23551_/B vssd1 vssd1 vccd1 vccd1 _23552_/A sky130_fd_sc_hd__and2_1
X_20763_ _20763_/A vssd1 vssd1 vccd1 vccd1 _20763_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_925 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22502_ _22502_/A vssd1 vssd1 vccd1 vccd1 _22502_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_26270_ _20257_/X _26270_/D vssd1 vssd1 vccd1 vccd1 _26270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23482_ _23482_/A vssd1 vssd1 vccd1 vccd1 _23482_/X sky130_fd_sc_hd__clkbuf_2
X_20694_ _20684_/X _20685_/X _20686_/X _20687_/X _20689_/X _20691_/X vssd1 vssd1 vccd1
+ vccd1 _20695_/A sky130_fd_sc_hd__mux4_1
X_25221_ _25221_/A _25221_/B vssd1 vssd1 vccd1 vccd1 _25221_/Y sky130_fd_sc_hd__nand2_1
X_22433_ _22433_/A vssd1 vssd1 vccd1 vccd1 _22433_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25152_ _27694_/Q _25142_/X _25151_/Y _25132_/X vssd1 vssd1 vccd1 vccd1 _27694_/D
+ sky130_fd_sc_hd__o211a_1
X_22364_ _22364_/A vssd1 vssd1 vccd1 vccd1 _22364_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24103_ _24103_/A vssd1 vssd1 vccd1 vccd1 _27326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21315_ _21301_/X _21302_/X _21303_/X _21304_/X _21307_/X _21310_/X vssd1 vssd1 vccd1
+ vccd1 _21316_/A sky130_fd_sc_hd__mux4_1
X_25083_ _27975_/A _25082_/X _25104_/S vssd1 vssd1 vccd1 vccd1 _25084_/A sky130_fd_sc_hd__mux2_1
X_22295_ _22280_/X _22282_/X _22284_/X _22286_/X _22287_/X _22288_/X vssd1 vssd1 vccd1
+ vccd1 _22296_/A sky130_fd_sc_hd__mux4_1
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24034_ _27095_/Q _24001_/X _24002_/X _27127_/Q _24003_/X vssd1 vssd1 vccd1 vccd1
+ _24034_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21246_ _21246_/A vssd1 vssd1 vccd1 vccd1 _21246_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21177_ _21163_/X _21164_/X _21165_/X _21166_/X _21167_/X _21168_/X vssd1 vssd1 vccd1
+ vccd1 _21178_/A sky130_fd_sc_hd__mux4_1
XFILLER_85_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20128_ _20114_/X _20115_/X _20116_/X _20117_/X _20118_/X _20119_/X vssd1 vssd1 vccd1
+ vccd1 _20129_/A sky130_fd_sc_hd__mux4_1
X_25985_ _25985_/CLK _25985_/D vssd1 vssd1 vccd1 vccd1 _25985_/Q sky130_fd_sc_hd__dfxtp_1
X_12950_ _27820_/Q _12952_/B vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__and2_1
XFILLER_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27724_ _27750_/CLK _27724_/D vssd1 vssd1 vccd1 vccd1 _27724_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ _20059_/A vssd1 vssd1 vccd1 vccd1 _20059_/X sky130_fd_sc_hd__clkbuf_1
X_24936_ _25580_/A _24941_/C vssd1 vssd1 vccd1 vccd1 _24937_/B sky130_fd_sc_hd__xnor2_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27655_ _27658_/CLK _27655_/D vssd1 vssd1 vccd1 vccd1 _27655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24867_ _27763_/Q _27762_/Q _24867_/C vssd1 vssd1 vccd1 vccd1 _24873_/B sky130_fd_sc_hd__and3_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _14497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _14511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26606_ _21436_/X _26606_/D vssd1 vssd1 vccd1 vccd1 _26606_/Q sky130_fd_sc_hd__dfxtp_1
X_14620_ _15781_/A _14620_/B vssd1 vssd1 vccd1 vccd1 _14620_/Y sky130_fd_sc_hd__nor2_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _14801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_234 _17321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_23818_ _27832_/Q _27136_/Q _25881_/Q _25849_/Q _23777_/X _23802_/X vssd1 vssd1 vccd1
+ vccd1 _23818_/X sky130_fd_sc_hd__mux4_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 _27423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_24798_ _24861_/A vssd1 vssd1 vccd1 vccd1 _24798_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27586_ _27587_/CLK _27586_/D vssd1 vssd1 vccd1 vccd1 _27586_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _26815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_763 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14551_ _26613_/Q _14549_/X _14536_/X _14550_/Y vssd1 vssd1 vccd1 vccd1 _26613_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA_267 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23749_ _23929_/A vssd1 vssd1 vccd1 vccd1 _23749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_278 input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_26537_ _21190_/X _26537_/D vssd1 vssd1 vccd1 vccd1 _26537_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _14471_/A vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14482_ _14482_/A vssd1 vssd1 vccd1 vccd1 _15745_/A sky130_fd_sc_hd__buf_2
X_17270_ _17242_/X _17269_/X _17220_/X vssd1 vssd1 vccd1 vccd1 _17270_/X sky130_fd_sc_hd__a21bo_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26468_ _20950_/X _26468_/D vssd1 vssd1 vccd1 vccd1 _26468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13433_ _13857_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13433_/Y sky130_fd_sc_hd__nor2_1
X_16221_ _26047_/Q _16221_/B _16221_/C vssd1 vssd1 vccd1 vccd1 _16221_/X sky130_fd_sc_hd__and3_1
X_25419_ _25419_/A vssd1 vssd1 vccd1 vccd1 _27747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26399_ _20701_/X _26399_/D vssd1 vssd1 vccd1 vccd1 _26399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ _26064_/Q vssd1 vssd1 vccd1 vccd1 _16152_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ _26988_/Q _13363_/X _13367_/S vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15103_ _15103_/A vssd1 vssd1 vccd1 vccd1 _15112_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_182_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16083_ _16625_/B vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13295_ _13295_/A vssd1 vssd1 vccd1 vccd1 _27013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15034_ _15771_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15034_/Y sky130_fd_sc_hd__nor2_1
X_19911_ _19911_/A vssd1 vssd1 vccd1 vccd1 _19911_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19842_ _19831_/X _19833_/X _19835_/X _19837_/X _19838_/X _19839_/X vssd1 vssd1 vccd1
+ vccd1 _19843_/A sky130_fd_sc_hd__mux4_1
XFILLER_69_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19773_ _19773_/A vssd1 vssd1 vccd1 vccd1 _19773_/X sky130_fd_sc_hd__clkbuf_1
X_16985_ _17220_/A vssd1 vssd1 vccd1 vccd1 _16985_/X sky130_fd_sc_hd__clkbuf_2
X_18724_ _26024_/Q _17721_/X _18724_/S vssd1 vssd1 vccd1 vccd1 _18725_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_1164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15936_ _15937_/A vssd1 vssd1 vccd1 vccd1 _15936_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18655_ _25993_/Q _17724_/X _18663_/S vssd1 vssd1 vccd1 vccd1 _18656_/A sky130_fd_sc_hd__mux2_1
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15867_ _15868_/A vssd1 vssd1 vccd1 vccd1 _15867_/Y sky130_fd_sc_hd__inv_2
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17606_ _17428_/X _25876_/Q _17612_/S vssd1 vssd1 vccd1 vccd1 _17607_/A sky130_fd_sc_hd__mux2_1
X_14818_ _26520_/Q _13325_/X _14824_/S vssd1 vssd1 vccd1 vccd1 _14819_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ _24640_/A _18601_/A vssd1 vssd1 vccd1 vccd1 _18605_/A sky130_fd_sc_hd__or2_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _15798_/A vssd1 vssd1 vccd1 vccd1 _26100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17537_ _17537_/A vssd1 vssd1 vccd1 vccd1 _25845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14749_ _14749_/A vssd1 vssd1 vccd1 vccd1 _26542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17468_ _17468_/A vssd1 vssd1 vccd1 vccd1 _25824_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19207_ _19158_/X _19206_/X _19089_/X vssd1 vssd1 vccd1 vccd1 _19207_/X sky130_fd_sc_hd__o21a_1
X_16419_ _16710_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16433_/A sky130_fd_sc_hd__or2_1
Xrepeater81 _27427_/CLK vssd1 vssd1 vccd1 vccd1 _27088_/CLK sky130_fd_sc_hd__clkbuf_1
Xrepeater92 _26001_/CLK vssd1 vssd1 vccd1 vccd1 _25895_/CLK sky130_fd_sc_hd__clkbuf_1
X_17399_ _20800_/A vssd1 vssd1 vccd1 vccd1 _25659_/A sky130_fd_sc_hd__buf_6
X_19138_ _18929_/X _19137_/X _18932_/X vssd1 vssd1 vccd1 vccd1 _19138_/X sky130_fd_sc_hd__o21a_1
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19069_ _18895_/X _19064_/X _19066_/X _19068_/X _19023_/X vssd1 vssd1 vccd1 vccd1
+ _19083_/B sky130_fd_sc_hd__a221o_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21100_ _21100_/A vssd1 vssd1 vccd1 vccd1 _21100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_22080_ _22080_/A vssd1 vssd1 vccd1 vccd1 _22080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21031_ _21023_/X _21024_/X _21025_/X _21026_/X _21027_/X _21028_/X vssd1 vssd1 vccd1
+ vccd1 _21032_/A sky130_fd_sc_hd__mux4_1
XFILLER_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25770_ _25792_/A vssd1 vssd1 vccd1 vccd1 _25779_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22982_ _23030_/A vssd1 vssd1 vccd1 vccd1 _22982_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21933_ _22019_/A vssd1 vssd1 vccd1 vccd1 _21999_/A sky130_fd_sc_hd__clkbuf_2
X_24721_ _27189_/Q _24725_/B vssd1 vssd1 vccd1 vccd1 _24721_/X sky130_fd_sc_hd__or2_1
XFILLER_41_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24652_ _27163_/Q _24658_/B vssd1 vssd1 vccd1 vccd1 _24652_/X sky130_fd_sc_hd__or2_1
X_27440_ _27443_/CLK _27440_/D vssd1 vssd1 vccd1 vccd1 _27440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21864_ _21912_/A vssd1 vssd1 vccd1 vccd1 _21864_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23603_ _23603_/A vssd1 vssd1 vccd1 vccd1 _27220_/D sky130_fd_sc_hd__clkbuf_1
X_20815_ _20815_/A vssd1 vssd1 vccd1 vccd1 _20815_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24583_ _27652_/Q _24587_/B vssd1 vssd1 vccd1 vccd1 _24584_/A sky130_fd_sc_hd__and2_1
X_27371_ _27480_/CLK _27371_/D vssd1 vssd1 vccd1 vccd1 _27371_/Q sky130_fd_sc_hd__dfxtp_1
X_21795_ _21827_/A vssd1 vssd1 vccd1 vccd1 _21795_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_430 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26322_ _20439_/X _26322_/D vssd1 vssd1 vccd1 vccd1 _26322_/Q sky130_fd_sc_hd__dfxtp_1
X_23534_ _23543_/A _23534_/B vssd1 vssd1 vccd1 vccd1 _23535_/A sky130_fd_sc_hd__and2_1
XFILLER_196_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20746_ _20738_/X _20739_/X _20740_/X _20741_/X _20742_/X _20743_/X vssd1 vssd1 vccd1
+ vccd1 _20747_/A sky130_fd_sc_hd__mux4_1
XFILLER_169_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26253_ _20197_/X _26253_/D vssd1 vssd1 vccd1 vccd1 _26253_/Q sky130_fd_sc_hd__dfxtp_1
X_23465_ _27179_/Q _23470_/B vssd1 vssd1 vccd1 vccd1 _23465_/X sky130_fd_sc_hd__or2_1
XFILLER_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20677_ _20677_/A vssd1 vssd1 vccd1 vccd1 _20677_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25204_ _25198_/A _25197_/B _25197_/A vssd1 vssd1 vccd1 vccd1 _25205_/B sky130_fd_sc_hd__a21boi_1
X_22416_ _22416_/A vssd1 vssd1 vccd1 vccd1 _22416_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26184_ _19955_/X _26184_/D vssd1 vssd1 vccd1 vccd1 _26184_/Q sky130_fd_sc_hd__dfxtp_1
X_23396_ _24776_/A _27249_/Q _23394_/Y _27777_/Q _23395_/X vssd1 vssd1 vccd1 vccd1
+ _23409_/A sky130_fd_sc_hd__a221o_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_546 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25135_ _27523_/Q _27491_/Q vssd1 vssd1 vccd1 vccd1 _25149_/A sky130_fd_sc_hd__or2_1
X_22347_ _22347_/A vssd1 vssd1 vccd1 vccd1 _22347_/X sky130_fd_sc_hd__clkbuf_1
X_27957__443 vssd1 vssd1 vccd1 vccd1 _27957__443/HI _27957_/A sky130_fd_sc_hd__conb_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25066_ _25064_/X _25065_/X _25074_/S vssd1 vssd1 vccd1 vccd1 _25066_/X sky130_fd_sc_hd__mux2_1
X_13080_ _13080_/A vssd1 vssd1 vccd1 vccd1 _27061_/D sky130_fd_sc_hd__clkbuf_1
X_22278_ _22278_/A vssd1 vssd1 vccd1 vccd1 _22278_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24017_ _24015_/X _24016_/X _24031_/S vssd1 vssd1 vccd1 vccd1 _24017_/X sky130_fd_sc_hd__mux2_1
X_21229_ _22537_/A vssd1 vssd1 vccd1 vccd1 _21579_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16770_ _16778_/A _16778_/B vssd1 vssd1 vccd1 vccd1 _16770_/Y sky130_fd_sc_hd__xnor2_1
X_13982_ _26800_/Q _13969_/X _13965_/X _13981_/Y vssd1 vssd1 vccd1 vccd1 _26800_/D
+ sky130_fd_sc_hd__a31o_1
X_25968_ _26059_/CLK _25968_/D vssd1 vssd1 vccd1 vccd1 _25968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15721_ _24980_/S vssd1 vssd1 vccd1 vccd1 _15721_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27707_ _27709_/CLK _27707_/D vssd1 vssd1 vccd1 vccd1 _27707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24919_ _24925_/C _24919_/B vssd1 vssd1 vccd1 vccd1 _24920_/B sky130_fd_sc_hd__or2_1
X_12933_ input20/X _27858_/Q _12933_/S vssd1 vssd1 vccd1 vccd1 _12934_/B sky130_fd_sc_hd__mux2_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_25899_ _27154_/CLK _25899_/D vssd1 vssd1 vccd1 vccd1 _25899_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _26546_/Q _26514_/Q _26482_/Q _27058_/Q _18392_/X _18418_/X vssd1 vssd1 vccd1
+ vccd1 _18440_/X sky130_fd_sc_hd__mux4_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27638_ _27720_/CLK _27638_/D vssd1 vssd1 vccd1 vccd1 _27638_/Q sky130_fd_sc_hd__dfxtp_1
X_15652_ _13128_/X _26157_/Q _15656_/S vssd1 vssd1 vccd1 vccd1 _15653_/A sky130_fd_sc_hd__mux2_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _15764_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14603_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _17827_/X _18370_/X _17838_/X vssd1 vssd1 vccd1 vccd1 _18371_/X sky130_fd_sc_hd__o21a_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15583_ _15583_/A vssd1 vssd1 vccd1 vccd1 _26188_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27569_ _27569_/CLK _27569_/D vssd1 vssd1 vccd1 vccd1 _27569_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _25358_/B vssd1 vssd1 vccd1 vccd1 _17367_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_109_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14534_ _15695_/D _14534_/B vssd1 vssd1 vccd1 vccd1 _14552_/A sky130_fd_sc_hd__nand2b_2
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17253_ _27846_/Q _27150_/Q _25895_/Q _25863_/Q _17203_/X _17252_/X vssd1 vssd1 vccd1
+ vccd1 _17253_/X sky130_fd_sc_hd__mux4_1
XFILLER_144_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14465_ _15732_/A _14465_/B vssd1 vssd1 vccd1 vccd1 _14465_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ _23035_/A _16233_/B vssd1 vssd1 vccd1 vccd1 _16204_/Y sky130_fd_sc_hd__nor2_1
X_13416_ _13416_/A vssd1 vssd1 vccd1 vccd1 _26972_/D sky130_fd_sc_hd__clkbuf_1
X_14396_ _14396_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14396_/Y sky130_fd_sc_hd__nor2_1
X_17184_ _17177_/X _17178_/X _17180_/X _17183_/X vssd1 vssd1 vccd1 vccd1 _17184_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16135_ _16131_/X _16133_/Y _16134_/X _16266_/A vssd1 vssd1 vccd1 vccd1 _16593_/B
+ sky130_fd_sc_hd__a31o_1
X_13347_ _14737_/A vssd1 vssd1 vccd1 vccd1 _13347_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13278_ _27020_/Q _13133_/X _13280_/S vssd1 vssd1 vccd1 vccd1 _13279_/A sky130_fd_sc_hd__mux2_1
X_16066_ _16066_/A _16066_/B _16066_/C vssd1 vssd1 vccd1 vccd1 _16457_/B sky130_fd_sc_hd__and3_1
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15017_ _15754_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _15017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19825_ _19825_/A vssd1 vssd1 vccd1 vccd1 _19825_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19756_ _19745_/X _19747_/X _19749_/X _19751_/X _19752_/X _19753_/X vssd1 vssd1 vccd1
+ vccd1 _19757_/A sky130_fd_sc_hd__mux4_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16968_ _27592_/Q vssd1 vssd1 vccd1 vccd1 _16979_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18707_ _26016_/Q _17696_/X _18713_/S vssd1 vssd1 vccd1 vccd1 _18708_/A sky130_fd_sc_hd__mux2_1
X_15919_ _15925_/A vssd1 vssd1 vccd1 vccd1 _15924_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19687_ _19687_/A vssd1 vssd1 vccd1 vccd1 _19687_/X sky130_fd_sc_hd__clkbuf_1
X_16899_ _16077_/X _16308_/A _16790_/B _16087_/X vssd1 vssd1 vccd1 vccd1 _16899_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18638_ _18638_/A vssd1 vssd1 vccd1 vccd1 _25985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18569_ _26841_/Q _26809_/Q _26777_/Q _26745_/Q _17832_/X _17835_/X vssd1 vssd1 vccd1
+ vccd1 _18569_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20600_ _20600_/A vssd1 vssd1 vccd1 vccd1 _20600_/X sky130_fd_sc_hd__clkbuf_1
X_21580_ _21647_/A vssd1 vssd1 vccd1 vccd1 _21580_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20531_ _20598_/A vssd1 vssd1 vccd1 vccd1 _20531_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23250_ _17520_/X _27160_/Q _23252_/S vssd1 vssd1 vccd1 vccd1 _23251_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20462_ _20445_/X _20447_/X _20449_/X _20451_/X _20452_/X _20453_/X vssd1 vssd1 vccd1
+ vccd1 _20463_/A sky130_fd_sc_hd__mux4_1
XFILLER_193_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22201_ _22249_/A vssd1 vssd1 vccd1 vccd1 _22201_/X sky130_fd_sc_hd__clkbuf_2
X_23181_ _23181_/A vssd1 vssd1 vccd1 vccd1 _27129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20393_ _20425_/A vssd1 vssd1 vccd1 vccd1 _20393_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22132_ _22132_/A vssd1 vssd1 vccd1 vccd1 _22132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22063_ _22051_/X _22052_/X _22053_/X _22054_/X _22055_/X _22056_/X vssd1 vssd1 vccd1
+ vccd1 _22064_/A sky130_fd_sc_hd__mux4_1
X_26940_ _22600_/X _26940_/D vssd1 vssd1 vccd1 vccd1 _26940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21014_ _21014_/A vssd1 vssd1 vccd1 vccd1 _21014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_26871_ _22358_/X _26871_/D vssd1 vssd1 vccd1 vccd1 _26871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25822_ _27077_/CLK _25822_/D vssd1 vssd1 vccd1 vccd1 _25822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22965_ _22955_/X _22956_/X _22957_/X _22958_/X _22960_/X _22962_/X vssd1 vssd1 vccd1
+ vccd1 _22966_/A sky130_fd_sc_hd__mux4_1
X_25753_ _17447_/X _27833_/Q _25757_/S vssd1 vssd1 vccd1 vccd1 _25754_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_24704_ _24398_/A _24700_/X _24702_/X _24703_/X vssd1 vssd1 vccd1 vccd1 _27598_/D
+ sky130_fd_sc_hd__o211a_1
X_21916_ _21985_/A vssd1 vssd1 vccd1 vccd1 _21916_/X sky130_fd_sc_hd__clkbuf_2
X_25684_ _25684_/A vssd1 vssd1 vccd1 vccd1 _25684_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22896_ _22944_/A vssd1 vssd1 vccd1 vccd1 _22896_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_27423_ _27423_/CLK _27423_/D vssd1 vssd1 vccd1 vccd1 _27423_/Q sky130_fd_sc_hd__dfxtp_1
X_21847_ _22019_/A vssd1 vssd1 vccd1 vccd1 _21913_/A sky130_fd_sc_hd__buf_2
X_24635_ _24635_/A _24635_/B vssd1 vssd1 vccd1 vccd1 _24636_/C sky130_fd_sc_hd__nand2_1
XFILLER_167_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24566_ _24566_/A vssd1 vssd1 vccd1 vccd1 _27544_/D sky130_fd_sc_hd__clkbuf_1
X_27354_ _27447_/CLK _27354_/D vssd1 vssd1 vccd1 vccd1 _27354_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21778_ _21826_/A vssd1 vssd1 vccd1 vccd1 _21778_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26305_ _20383_/X _26305_/D vssd1 vssd1 vccd1 vccd1 _26305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20729_ _20729_/A vssd1 vssd1 vccd1 vccd1 _20729_/X sky130_fd_sc_hd__clkbuf_1
X_23517_ _24831_/B _27197_/Q _23525_/S vssd1 vssd1 vccd1 vccd1 _23518_/B sky130_fd_sc_hd__mux2_1
X_27285_ _27285_/CLK _27285_/D vssd1 vssd1 vccd1 vccd1 _27285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24497_ _24522_/A vssd1 vssd1 vccd1 vccd1 _24633_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_184_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14257_/A vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23448_ input10/X _23442_/X _23446_/X _23447_/X vssd1 vssd1 vccd1 vccd1 _27172_/D
+ sky130_fd_sc_hd__o211a_1
X_26236_ _20139_/X _26236_/D vssd1 vssd1 vccd1 vccd1 _26236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13201_ _27277_/Q _13201_/B vssd1 vssd1 vccd1 vccd1 _13201_/X sky130_fd_sc_hd__and2_1
XFILLER_137_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14181_ _14220_/A vssd1 vssd1 vccd1 vccd1 _14181_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23379_ _24877_/A vssd1 vssd1 vccd1 vccd1 _24765_/A sky130_fd_sc_hd__clkinv_2
X_26167_ _19893_/X _26167_/D vssd1 vssd1 vccd1 vccd1 _26167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ _27353_/Q _13529_/A _13530_/A _27321_/Q _13131_/X vssd1 vssd1 vccd1 vccd1
+ _14753_/A sky130_fd_sc_hd__a221o_4
XFILLER_174_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_25118_ _27540_/Q _27519_/Q _18612_/B _18610_/X vssd1 vssd1 vccd1 vccd1 _25122_/A
+ sky130_fd_sc_hd__a31o_1
X_26098_ _19655_/X _26098_/D vssd1 vssd1 vccd1 vccd1 _26098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17940_ _18483_/A vssd1 vssd1 vccd1 vccd1 _17940_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25049_ _27971_/A _25048_/X _25067_/S vssd1 vssd1 vccd1 vccd1 _25050_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13063_ _13063_/A vssd1 vssd1 vccd1 vccd1 _13063_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_152_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17871_ _26139_/Q _26075_/Q _27003_/Q _26971_/Q _17870_/X _17824_/X vssd1 vssd1 vccd1
+ vccd1 _17872_/A sky130_fd_sc_hd__mux4_1
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19610_ _19626_/A vssd1 vssd1 vccd1 vccd1 _19610_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16822_ _16822_/A _16801_/A vssd1 vssd1 vccd1 vccd1 _16822_/X sky130_fd_sc_hd__or2b_1
XFILLER_78_477 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19541_ _26168_/Q _26104_/Q _27032_/Q _27000_/Q _19460_/X _19482_/X vssd1 vssd1 vccd1
+ vccd1 _19542_/B sky130_fd_sc_hd__mux4_1
X_16753_ _16753_/A _16753_/B _16755_/A vssd1 vssd1 vccd1 vccd1 _16753_/X sky130_fd_sc_hd__or3b_1
X_13965_ _14038_/A vssd1 vssd1 vccd1 vccd1 _13965_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15704_ _26135_/Q _15040_/X _15697_/X _15703_/Y vssd1 vssd1 vccd1 vccd1 _26135_/D
+ sky130_fd_sc_hd__a31o_1
X_19472_ _19472_/A vssd1 vssd1 vccd1 vccd1 _26068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16684_ _16481_/A _16606_/Y _16450_/A _16450_/B vssd1 vssd1 vccd1 vccd1 _16684_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_13896_ _26828_/Q _13893_/X _13886_/X _13895_/Y vssd1 vssd1 vccd1 vccd1 _26828_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18423_ _18509_/A _18423_/B _18423_/C vssd1 vssd1 vccd1 vccd1 _18424_/A sky130_fd_sc_hd__and3_1
XFILLER_59_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ _15635_/A vssd1 vssd1 vccd1 vccd1 _26165_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _18354_/A vssd1 vssd1 vccd1 vccd1 _25964_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15566_ _15566_/A vssd1 vssd1 vccd1 vccd1 _26196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17303_/X _17304_/X _17281_/X vssd1 vssd1 vccd1 vccd1 _17305_/X sky130_fd_sc_hd__a21bo_1
XFILLER_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14517_ _26623_/Q _14514_/X _14510_/X _14516_/Y vssd1 vssd1 vccd1 vccd1 _26623_/D
+ sky130_fd_sc_hd__a31o_1
X_18285_ _18285_/A vssd1 vssd1 vccd1 vccd1 _18285_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15497_ _13099_/X _26226_/Q _15501_/S vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__mux2_1
X_17236_ _27213_/Q _17235_/X _17250_/S vssd1 vssd1 vccd1 vccd1 _17237_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14448_ _14448_/A vssd1 vssd1 vccd1 vccd1 _15723_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17167_ _25925_/Q _25991_/Q _17193_/S vssd1 vssd1 vccd1 vccd1 _17168_/B sky130_fd_sc_hd__mux2_1
X_14379_ _14441_/A vssd1 vssd1 vccd1 vccd1 _14379_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16118_ _16274_/B _16274_/C vssd1 vssd1 vccd1 vccd1 _16119_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17098_ _17220_/A vssd1 vssd1 vccd1 vccd1 _17098_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16049_ _27478_/Q _27374_/Q vssd1 vssd1 vccd1 vccd1 _16049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19808_ _19796_/X _19797_/X _19798_/X _19799_/X _19800_/X _19801_/X vssd1 vssd1 vccd1
+ vccd1 _19809_/A sky130_fd_sc_hd__mux4_1
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19739_ _19739_/A vssd1 vssd1 vccd1 vccd1 _19739_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22750_ _22750_/A vssd1 vssd1 vccd1 vccd1 _22750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21701_ _21689_/X _21690_/X _21691_/X _21692_/X _21693_/X _21694_/X vssd1 vssd1 vccd1
+ vccd1 _21702_/A sky130_fd_sc_hd__mux4_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22681_ _22697_/A vssd1 vssd1 vccd1 vccd1 _22681_/X sky130_fd_sc_hd__clkbuf_1
X_24420_ _27610_/Q _24422_/B vssd1 vssd1 vccd1 vccd1 _24421_/A sky130_fd_sc_hd__and2_1
X_21632_ _21648_/A vssd1 vssd1 vccd1 vccd1 _21632_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24351_ _24351_/A vssd1 vssd1 vccd1 vccd1 _27458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21563_ _21563_/A vssd1 vssd1 vccd1 vccd1 _21563_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23302_ _27751_/Q vssd1 vssd1 vccd1 vccd1 _23302_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20514_ _20514_/A vssd1 vssd1 vccd1 vccd1 _20514_/X sky130_fd_sc_hd__clkbuf_1
X_27070_ _27413_/CLK _27070_/D vssd1 vssd1 vccd1 vccd1 _27070_/Q sky130_fd_sc_hd__dfxtp_1
X_24282_ _16166_/X _16168_/Y _16169_/X _24279_/X vssd1 vssd1 vccd1 vccd1 _27418_/D
+ sky130_fd_sc_hd__o31a_1
X_21494_ _21561_/A vssd1 vssd1 vccd1 vccd1 _21494_/X sky130_fd_sc_hd__clkbuf_1
X_23233_ _17495_/X _27152_/Q _23237_/S vssd1 vssd1 vccd1 vccd1 _23234_/A sky130_fd_sc_hd__mux2_1
X_26021_ _27077_/CLK _26021_/D vssd1 vssd1 vccd1 vccd1 _26021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20445_ _20512_/A vssd1 vssd1 vccd1 vccd1 _20445_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_23164_ _23164_/A vssd1 vssd1 vccd1 vccd1 _27121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20376_ _20424_/A vssd1 vssd1 vccd1 vccd1 _20376_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22115_ _22103_/X _22106_/X _22109_/X _22112_/X _22113_/X _22114_/X vssd1 vssd1 vccd1
+ vccd1 _22116_/A sky130_fd_sc_hd__mux4_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23095_ _27091_/Q _17756_/X _23103_/S vssd1 vssd1 vccd1 vccd1 _23096_/A sky130_fd_sc_hd__mux2_1
X_27972_ _27972_/A _15939_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
XFILLER_133_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22046_ _22046_/A vssd1 vssd1 vccd1 vccd1 _22046_/X sky130_fd_sc_hd__clkbuf_1
X_26923_ _22534_/X _26923_/D vssd1 vssd1 vccd1 vccd1 _26923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_657 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_26854_ _22298_/X _26854_/D vssd1 vssd1 vccd1 vccd1 _26854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_436 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_25805_ _17523_/X _27857_/Q _25805_/S vssd1 vssd1 vccd1 vccd1 _25806_/A sky130_fd_sc_hd__mux2_1
X_26785_ _22058_/X _26785_/D vssd1 vssd1 vccd1 vccd1 _26785_/Q sky130_fd_sc_hd__dfxtp_1
X_23997_ _23997_/A vssd1 vssd1 vccd1 vccd1 _24032_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13750_ _13778_/A vssd1 vssd1 vccd1 vccd1 _13750_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_25736_ _25792_/A vssd1 vssd1 vccd1 vccd1 _25805_/S sky130_fd_sc_hd__buf_2
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22948_ _22948_/A vssd1 vssd1 vccd1 vccd1 _22948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_828 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13681_ _26904_/Q _13665_/X _13676_/X _13680_/Y vssd1 vssd1 vccd1 vccd1 _26904_/D
+ sky130_fd_sc_hd__a31o_1
X_25667_ _25654_/X _25656_/X _25658_/X _25660_/X _25661_/X _25662_/X vssd1 vssd1 vccd1
+ vccd1 _25668_/A sky130_fd_sc_hd__mux4_1
X_22879_ _22869_/X _22870_/X _22871_/X _22872_/X _22874_/X _22876_/X vssd1 vssd1 vccd1
+ vccd1 _22880_/A sky130_fd_sc_hd__mux4_1
XFILLER_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27406_ _27406_/CLK _27406_/D vssd1 vssd1 vccd1 vccd1 _27406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15420_ _15477_/S vssd1 vssd1 vccd1 vccd1 _15429_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24618_ _27668_/Q _24620_/B vssd1 vssd1 vccd1 vccd1 _24619_/A sky130_fd_sc_hd__and2_1
XFILLER_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25598_ _24267_/A _25440_/X _25442_/X _24957_/B _24384_/A vssd1 vssd1 vccd1 vccd1
+ _25598_/X sky130_fd_sc_hd__o311a_1
XFILLER_169_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15351_ _14731_/X _26291_/Q _15357_/S vssd1 vssd1 vccd1 vccd1 _15352_/A sky130_fd_sc_hd__mux2_1
X_27337_ _27338_/CLK _27337_/D vssd1 vssd1 vccd1 vccd1 _27337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_24549_ _24552_/A _24549_/B vssd1 vssd1 vccd1 vccd1 _24550_/A sky130_fd_sc_hd__and2_1
XFILLER_184_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14302_ _14390_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14302_/Y sky130_fd_sc_hd__nor2_1
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18070_ _18483_/A vssd1 vssd1 vccd1 vccd1 _18070_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ _26321_/Q _13347_/X _15284_/S vssd1 vssd1 vccd1 vccd1 _15283_/A sky130_fd_sc_hd__mux2_1
X_27268_ _27480_/CLK _27268_/D vssd1 vssd1 vccd1 vccd1 _27268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17021_ _25812_/Q _26011_/Q _17061_/A vssd1 vssd1 vccd1 vccd1 _17021_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14233_ _26715_/Q _14225_/X _14158_/B _14232_/Y vssd1 vssd1 vccd1 vccd1 _26715_/D
+ sky130_fd_sc_hd__a31o_1
X_26219_ _20075_/X _26219_/D vssd1 vssd1 vccd1 vccd1 _26219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_27199_ _27207_/CLK _27199_/D vssd1 vssd1 vccd1 vccd1 _27199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _14342_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14164_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13115_ _27356_/Q _13090_/X _13091_/X _27324_/Q _13114_/X vssd1 vssd1 vccd1 vccd1
+ _14743_/A sky130_fd_sc_hd__a221o_2
X_14095_ _26767_/Q _14090_/X _14093_/X _14094_/Y vssd1 vssd1 vccd1 vccd1 _26767_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18972_ _19412_/A vssd1 vssd1 vccd1 vccd1 _18972_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17923_ _26941_/Q _26909_/Q _26877_/Q _26845_/Q _17922_/X _17791_/X vssd1 vssd1 vccd1
+ vccd1 _17923_/X sky130_fd_sc_hd__mux4_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _27266_/Q vssd1 vssd1 vccd1 vccd1 _13672_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17854_ _18285_/A vssd1 vssd1 vccd1 vccd1 _17854_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_1179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16805_ _16805_/A _16805_/B vssd1 vssd1 vccd1 vccd1 _16805_/Y sky130_fd_sc_hd__xnor2_1
X_17785_ _18481_/A vssd1 vssd1 vccd1 vccd1 _17785_/X sky130_fd_sc_hd__buf_2
XFILLER_94_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14997_ _15736_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _14997_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_650 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19524_ _19524_/A _19524_/B vssd1 vssd1 vccd1 vccd1 _19524_/X sky130_fd_sc_hd__or2_1
X_16736_ _16738_/A _16732_/Y _16735_/X _16626_/A vssd1 vssd1 vccd1 vccd1 _24228_/A
+ sky130_fd_sc_hd__a22o_1
X_13948_ _26809_/Q _13933_/X _13944_/X _13947_/Y vssd1 vssd1 vccd1 vccd1 _26809_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_631 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19455_ _19431_/X _19454_/X _19387_/X vssd1 vssd1 vccd1 vccd1 _19455_/X sky130_fd_sc_hd__o21a_1
X_16667_ _16621_/X _16665_/X _16666_/Y vssd1 vssd1 vccd1 vccd1 _16667_/X sky130_fd_sc_hd__o21ba_1
X_13879_ _26834_/Q _13865_/X _13873_/X _13878_/Y vssd1 vssd1 vccd1 vccd1 _26834_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18406_ _18402_/X _18404_/X _18532_/S vssd1 vssd1 vccd1 vccd1 _18406_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15618_ _15618_/A vssd1 vssd1 vccd1 vccd1 _26172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_195_809 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19386_ _26705_/Q _26673_/Q _26641_/Q _26609_/Q _19317_/X _19385_/X vssd1 vssd1 vccd1
+ vccd1 _19386_/X sky130_fd_sc_hd__mux4_2
X_16598_ _16598_/A _16598_/B vssd1 vssd1 vccd1 vccd1 _16902_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18337_ _26830_/Q _26798_/Q _26766_/Q _26734_/Q _18387_/A _17810_/X vssd1 vssd1 vccd1
+ vccd1 _18337_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15549_ _13240_/X _26202_/Q _15549_/S vssd1 vssd1 vccd1 vccd1 _15550_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18268_ _27810_/Q _26571_/Q _26443_/Q _26123_/Q _18242_/X _18267_/X vssd1 vssd1 vccd1
+ vccd1 _18268_/X sky130_fd_sc_hd__mux4_2
XFILLER_147_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17219_ _25828_/Q _26027_/Q _17219_/S vssd1 vssd1 vccd1 vccd1 _17219_/X sky130_fd_sc_hd__mux2_1
X_18199_ _18380_/A vssd1 vssd1 vccd1 vccd1 _18199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_622 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20230_ _20216_/X _20217_/X _20218_/X _20219_/X _20220_/X _20221_/X vssd1 vssd1 vccd1
+ vccd1 _20231_/A sky130_fd_sc_hd__mux4_1
XFILLER_196_1070 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20161_ _20161_/A vssd1 vssd1 vccd1 vccd1 _20161_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20092_ _20076_/X _20077_/X _20078_/X _20079_/X _20081_/X _20083_/X vssd1 vssd1 vccd1
+ vccd1 _20093_/A sky130_fd_sc_hd__mux4_1
XFILLER_58_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23920_ _24014_/A vssd1 vssd1 vccd1 vccd1 _23920_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_28014__480 vssd1 vssd1 vccd1 vccd1 _28014__480/HI _28014_/A sky130_fd_sc_hd__conb_1
XFILLER_97_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23851_ _27836_/Q _27140_/Q _25885_/Q _25853_/Q _23826_/X _23850_/X vssd1 vssd1 vccd1
+ vccd1 _23851_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22802_ _22869_/A vssd1 vssd1 vccd1 vccd1 _22802_/X sky130_fd_sc_hd__clkbuf_1
X_26570_ _21312_/X _26570_/D vssd1 vssd1 vccd1 vccd1 _26570_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20994_ _21042_/A vssd1 vssd1 vccd1 vccd1 _20994_/X sky130_fd_sc_hd__clkbuf_1
X_23782_ _23780_/X _23781_/X _23797_/S vssd1 vssd1 vccd1 vccd1 _23782_/X sky130_fd_sc_hd__mux2_1
X_25521_ _27704_/Q _25509_/X _25510_/X vssd1 vssd1 vccd1 vccd1 _25521_/Y sky130_fd_sc_hd__a21oi_1
X_22733_ _22716_/X _22718_/X _22720_/X _22722_/X _22723_/X _22724_/X vssd1 vssd1 vccd1
+ vccd1 _22734_/A sky130_fd_sc_hd__mux4_1
XFILLER_168_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22664_ _22664_/A vssd1 vssd1 vccd1 vccd1 _22664_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_25452_ _25543_/A vssd1 vssd1 vccd1 vccd1 _25452_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21615_ _21647_/A vssd1 vssd1 vccd1 vccd1 _21615_/X sky130_fd_sc_hd__clkbuf_1
X_24403_ _24403_/A _24411_/B vssd1 vssd1 vccd1 vccd1 _24404_/A sky130_fd_sc_hd__and2_1
XFILLER_185_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22595_ _22611_/A vssd1 vssd1 vccd1 vccd1 _22595_/X sky130_fd_sc_hd__clkbuf_1
X_25383_ _27731_/Q input42/X _25391_/S vssd1 vssd1 vccd1 vccd1 _25384_/A sky130_fd_sc_hd__mux2_1
X_27122_ _27122_/CLK _27122_/D vssd1 vssd1 vccd1 vccd1 _27122_/Q sky130_fd_sc_hd__dfxtp_1
X_21546_ _21562_/A vssd1 vssd1 vccd1 vccd1 _21546_/X sky130_fd_sc_hd__clkbuf_1
X_24334_ _24334_/A vssd1 vssd1 vccd1 vccd1 _27450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_24265_ _25572_/A vssd1 vssd1 vccd1 vccd1 _25517_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_27053_ _22990_/X _27053_/D vssd1 vssd1 vccd1 vccd1 _27053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21477_ _21477_/A vssd1 vssd1 vccd1 vccd1 _21477_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23216_ _23216_/A vssd1 vssd1 vccd1 vccd1 _27144_/D sky130_fd_sc_hd__clkbuf_1
X_26004_ _27125_/CLK _26004_/D vssd1 vssd1 vccd1 vccd1 _26004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20428_ _25639_/A vssd1 vssd1 vccd1 vccd1 _20774_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24196_ _24196_/A vssd1 vssd1 vccd1 vccd1 _27368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_23147_ _23147_/A vssd1 vssd1 vccd1 vccd1 _27113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20359_ _20706_/A vssd1 vssd1 vccd1 vccd1 _20426_/A sky130_fd_sc_hd__buf_2
XFILLER_49_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_933 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_27955_ _27955_/A _15917_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
X_23078_ _23078_/A vssd1 vssd1 vccd1 vccd1 _27083_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22029_ _22016_/X _22018_/X _22020_/X _22022_/X _22023_/X _22024_/X vssd1 vssd1 vccd1
+ vccd1 _22030_/A sky130_fd_sc_hd__mux4_1
X_26906_ _22480_/X _26906_/D vssd1 vssd1 vccd1 vccd1 _26906_/Q sky130_fd_sc_hd__dfxtp_1
X_14920_ _14942_/A vssd1 vssd1 vccd1 vccd1 _14929_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_26837_ _22240_/X _26837_/D vssd1 vssd1 vccd1 vccd1 _26837_/Q sky130_fd_sc_hd__dfxtp_1
X_14851_ _26505_/Q _13373_/X _14857_/S vssd1 vssd1 vccd1 vccd1 _14852_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _13895_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13802_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17570_ _17570_/A vssd1 vssd1 vccd1 vccd1 _25860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26768_ _21994_/X _26768_/D vssd1 vssd1 vccd1 vccd1 _26768_/Q sky130_fd_sc_hd__dfxtp_1
X_14782_ _16235_/A vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_1137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16521_ _27399_/Q _16557_/B _16384_/X _14737_/A vssd1 vssd1 vccd1 vccd1 _16521_/X
+ sky130_fd_sc_hd__a22o_1
X_13733_ _13913_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13733_/Y sky130_fd_sc_hd__nor2_1
X_25719_ _25705_/X _25706_/X _25707_/X _25708_/X _25709_/X _25710_/X vssd1 vssd1 vccd1
+ vccd1 _25720_/A sky130_fd_sc_hd__mux4_1
XFILLER_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_26699_ _21756_/X _26699_/D vssd1 vssd1 vccd1 vccd1 _26699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19240_ _19399_/A vssd1 vssd1 vccd1 vccd1 _19240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_472 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16452_ _27391_/Q _16094_/A _16098_/A _25959_/Q _16451_/Y vssd1 vssd1 vccd1 vccd1
+ _16768_/B sky130_fd_sc_hd__a221o_2
X_13664_ _26909_/Q _13653_/X _13656_/X _13663_/Y vssd1 vssd1 vccd1 vccd1 _26909_/D
+ sky130_fd_sc_hd__a31o_1
X_15403_ _14807_/X _26267_/Q _15405_/S vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__mux2_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ _26407_/Q _26375_/Q _26343_/Q _26311_/Q _19170_/X _19100_/X vssd1 vssd1 vccd1
+ vccd1 _19171_/X sky130_fd_sc_hd__mux4_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _16383_/A _16383_/B vssd1 vssd1 vccd1 vccd1 _16715_/C sky130_fd_sc_hd__nand2_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13595_ _13602_/A vssd1 vssd1 vccd1 vccd1 _13649_/A sky130_fd_sc_hd__clkbuf_2
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ _18238_/A vssd1 vssd1 vccd1 vccd1 _18122_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15334_ _15045_/B _15334_/B _15334_/C vssd1 vssd1 vccd1 vccd1 _15551_/B sky130_fd_sc_hd__nand3b_2
XFILLER_184_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053_ _18053_/A vssd1 vssd1 vccd1 vccd1 _25951_/D sky130_fd_sc_hd__clkbuf_1
X_15265_ _26329_/Q _13319_/X _15273_/S vssd1 vssd1 vccd1 vccd1 _15266_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_4 _21142_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _17307_/A vssd1 vssd1 vccd1 vccd1 _17047_/S sky130_fd_sc_hd__buf_2
X_14216_ _14394_/A _14226_/B vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15196_ _15196_/A vssd1 vssd1 vccd1 vccd1 _26360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14147_ _14412_/A _14147_/B vssd1 vssd1 vccd1 vccd1 _14147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14078_ _26773_/Q _14076_/X _14064_/X _14077_/Y vssd1 vssd1 vccd1 vccd1 _26773_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_113_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18955_ _19385_/A vssd1 vssd1 vccd1 vccd1 _18955_/X sky130_fd_sc_hd__buf_2
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17906_ _17924_/A vssd1 vssd1 vccd1 vccd1 _18522_/S sky130_fd_sc_hd__buf_4
X_13029_ _13029_/A vssd1 vssd1 vccd1 vccd1 _13530_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18886_ _18814_/X _18885_/X _18821_/X vssd1 vssd1 vccd1 vccd1 _18886_/X sky130_fd_sc_hd__o21a_1
XFILLER_121_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17837_ _27596_/Q vssd1 vssd1 vccd1 vccd1 _18014_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17768_ _17768_/A vssd1 vssd1 vccd1 vccd1 _25940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ _16719_/A _16719_/B _16719_/C vssd1 vssd1 vccd1 vccd1 _16719_/Y sky130_fd_sc_hd__nand3_1
X_19507_ _26294_/Q _26262_/Q _26230_/Q _26198_/Q _19441_/X _19486_/X vssd1 vssd1 vccd1
+ vccd1 _19507_/X sky130_fd_sc_hd__mux4_1
XFILLER_23_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17699_ _27415_/Q vssd1 vssd1 vccd1 vccd1 _17699_/X sky130_fd_sc_hd__clkbuf_2
X_19438_ _19438_/A vssd1 vssd1 vccd1 vccd1 _19524_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19369_ _19501_/A _19369_/B vssd1 vssd1 vccd1 vccd1 _19369_/X sky130_fd_sc_hd__or2_1
XFILLER_50_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21400_ _21400_/A vssd1 vssd1 vccd1 vccd1 _21400_/X sky130_fd_sc_hd__clkbuf_1
X_22380_ _22380_/A vssd1 vssd1 vccd1 vccd1 _22380_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21331_ _21322_/X _21324_/X _21326_/X _21328_/X _21329_/X _21330_/X vssd1 vssd1 vccd1
+ vccd1 _21332_/A sky130_fd_sc_hd__mux4_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24050_ _27376_/Q _24050_/B vssd1 vssd1 vccd1 vccd1 _24051_/A sky130_fd_sc_hd__and2_1
XFILLER_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21262_ _21262_/A vssd1 vssd1 vccd1 vccd1 _21262_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_23001_ _22993_/X _22994_/X _22995_/X _22996_/X _22997_/X _22998_/X vssd1 vssd1 vccd1
+ vccd1 _23002_/A sky130_fd_sc_hd__mux4_1
XFILLER_132_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20213_ _20213_/A vssd1 vssd1 vccd1 vccd1 _20213_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21193_ _21179_/X _21180_/X _21181_/X _21182_/X _21183_/X _21184_/X vssd1 vssd1 vccd1
+ vccd1 _21194_/A sky130_fd_sc_hd__mux4_1
XFILLER_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20144_ _20130_/X _20131_/X _20132_/X _20133_/X _20134_/X _20135_/X vssd1 vssd1 vccd1
+ vccd1 _20145_/A sky130_fd_sc_hd__mux4_1
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_27740_ _27748_/CLK _27740_/D vssd1 vssd1 vccd1 vccd1 _27740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20075_ _20075_/A vssd1 vssd1 vccd1 vccd1 _20075_/X sky130_fd_sc_hd__clkbuf_1
X_24952_ _24962_/A _24952_/B vssd1 vssd1 vccd1 vccd1 _24952_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23903_ _23997_/A vssd1 vssd1 vccd1 vccd1 _23939_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_58_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_27671_ _27754_/CLK _27671_/D vssd1 vssd1 vccd1 vccd1 _27671_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_24883_ _24889_/A _24883_/B vssd1 vssd1 vccd1 vccd1 _24883_/Y sky130_fd_sc_hd__nand2_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater360 _25909_/CLK vssd1 vssd1 vccd1 vccd1 _27585_/CLK sky130_fd_sc_hd__clkbuf_1
X_26622_ _21488_/X _26622_/D vssd1 vssd1 vccd1 vccd1 _26622_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater371 _27682_/CLK vssd1 vssd1 vccd1 vccd1 _27224_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater382 _27450_/CLK vssd1 vssd1 vccd1 vccd1 _27352_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_23834_ _27834_/Q _27138_/Q _25883_/Q _25851_/Q _23826_/X _23802_/X vssd1 vssd1 vccd1
+ vccd1 _23834_/X sky130_fd_sc_hd__mux4_1
Xrepeater393 _27341_/CLK vssd1 vssd1 vccd1 vccd1 _27342_/CLK sky130_fd_sc_hd__clkbuf_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_26553_ _21250_/X _26553_/D vssd1 vssd1 vccd1 vccd1 _26553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _21149_/A vssd1 vssd1 vccd1 vccd1 _21042_/A sky130_fd_sc_hd__buf_2
X_23765_ _23862_/A vssd1 vssd1 vccd1 vccd1 _23765_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25504_ _25564_/A vssd1 vssd1 vccd1 vccd1 _25504_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22716_ _22783_/A vssd1 vssd1 vccd1 vccd1 _22716_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_26484_ _21006_/X _26484_/D vssd1 vssd1 vccd1 vccd1 _26484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_23696_ _23707_/A vssd1 vssd1 vccd1 vccd1 _23705_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25435_ _25569_/A vssd1 vssd1 vccd1 vccd1 _25435_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22647_ _22630_/X _22632_/X _22634_/X _22636_/X _22637_/X _22638_/X vssd1 vssd1 vccd1
+ vccd1 _22648_/A sky130_fd_sc_hd__mux4_1
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13380_ _26983_/Q _13379_/X _13383_/S vssd1 vssd1 vccd1 vccd1 _13381_/A sky130_fd_sc_hd__mux2_1
X_22578_ _22610_/A vssd1 vssd1 vccd1 vccd1 _22578_/X sky130_fd_sc_hd__clkbuf_1
X_25366_ _25366_/A vssd1 vssd1 vccd1 vccd1 _27723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27105_ _27105_/CLK _27105_/D vssd1 vssd1 vccd1 vccd1 _27105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_588 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_24317_ _27543_/Q _24317_/B vssd1 vssd1 vccd1 vccd1 _24318_/A sky130_fd_sc_hd__and2_1
X_21529_ _21561_/A vssd1 vssd1 vccd1 vccd1 _21529_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_25297_ _25297_/A vssd1 vssd1 vccd1 vccd1 _25297_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_27036_ _22932_/X _27036_/D vssd1 vssd1 vccd1 vccd1 _27036_/Q sky130_fd_sc_hd__dfxtp_1
X_15050_ _15050_/A vssd1 vssd1 vccd1 vccd1 _26425_/D sky130_fd_sc_hd__clkbuf_1
X_24248_ _24248_/A vssd1 vssd1 vccd1 vccd1 _27395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14001_ _14038_/A vssd1 vssd1 vccd1 vccd1 _14001_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_181_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_24179_ _24179_/A vssd1 vssd1 vccd1 vccd1 _27360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_433 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18740_ _26031_/Q _17744_/X _18746_/S vssd1 vssd1 vccd1 vccd1 _18741_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15952_ _15955_/A vssd1 vssd1 vccd1 vccd1 _15952_/Y sky130_fd_sc_hd__inv_2
X_27938_ _27938_/A _15945_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
XFILLER_163_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14903_ _14734_/X _26482_/Q _14907_/S vssd1 vssd1 vccd1 vccd1 _14904_/A sky130_fd_sc_hd__mux2_1
X_18671_ _18671_/A vssd1 vssd1 vccd1 vccd1 _26000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _15887_/A vssd1 vssd1 vccd1 vccd1 _15883_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _17622_/A vssd1 vssd1 vccd1 vccd1 _25883_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _14834_/A vssd1 vssd1 vccd1 vccd1 _26513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _17599_/S vssd1 vssd1 vccd1 vccd1 _17562_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_45_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14765_ _14765_/A vssd1 vssd1 vccd1 vccd1 _26537_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16504_ _16632_/B vssd1 vssd1 vccd1 vccd1 _16815_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _13897_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13716_/Y sky130_fd_sc_hd__nor2_1
X_17484_ _17484_/A vssd1 vssd1 vccd1 vccd1 _25829_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14696_ _15769_/A _14699_/B vssd1 vssd1 vccd1 vccd1 _14696_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19223_ _19223_/A vssd1 vssd1 vccd1 vccd1 _26057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_189_488 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16435_ _27389_/Q _16094_/X _16434_/X vssd1 vssd1 vccd1 vccd1 _16769_/B sky130_fd_sc_hd__a21oi_2
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _13917_/A _13647_/B vssd1 vssd1 vccd1 vccd1 _13647_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19154_ _19154_/A vssd1 vssd1 vccd1 vccd1 _26054_/D sky130_fd_sc_hd__clkbuf_1
X_16366_ _14515_/A _16400_/A _16067_/X _16364_/Y _16365_/Y vssd1 vssd1 vccd1 vccd1
+ _16745_/B sky130_fd_sc_hd__o221a_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _26939_/Q _13558_/X _13442_/B _13577_/Y vssd1 vssd1 vccd1 vccd1 _26939_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_185_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18105_ _26820_/Q _26788_/Q _26756_/Q _26724_/Q _18034_/X _18058_/X vssd1 vssd1 vccd1
+ vccd1 _18105_/X sky130_fd_sc_hd__mux4_1
X_15317_ _26305_/Q _13398_/X _15317_/S vssd1 vssd1 vccd1 vccd1 _15318_/A sky130_fd_sc_hd__mux2_1
X_19085_ _26820_/Q _26788_/Q _26756_/Q _26724_/Q _19039_/X _18967_/X vssd1 vssd1 vccd1
+ vccd1 _19086_/B sky130_fd_sc_hd__mux4_1
X_16297_ _27401_/Q _16297_/B vssd1 vssd1 vccd1 vccd1 _16297_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18036_ _18177_/A vssd1 vssd1 vccd1 vccd1 _18036_/X sky130_fd_sc_hd__buf_2
XFILLER_145_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15248_ _14791_/X _26336_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15249_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15179_ _15179_/A vssd1 vssd1 vccd1 vccd1 _26367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19987_ _19987_/A vssd1 vssd1 vccd1 vccd1 _19987_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18938_ _18969_/A _18938_/B vssd1 vssd1 vccd1 vccd1 _18938_/X sky130_fd_sc_hd__or2_1
.ends

