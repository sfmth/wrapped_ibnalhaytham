magic
tech sky130B
magscale 1 2
timestamp 1661612359
<< obsli1 >>
rect 1104 2159 111872 112625
<< obsm1 >>
rect 14 1504 112962 113280
<< metal2 >>
rect 1306 114354 1362 115154
rect 3238 114354 3294 115154
rect 5170 114354 5226 115154
rect 7102 114354 7158 115154
rect 9678 114354 9734 115154
rect 11610 114354 11666 115154
rect 13542 114354 13598 115154
rect 15474 114354 15530 115154
rect 18050 114354 18106 115154
rect 19982 114354 20038 115154
rect 21914 114354 21970 115154
rect 23846 114354 23902 115154
rect 26422 114354 26478 115154
rect 28354 114354 28410 115154
rect 30286 114354 30342 115154
rect 32218 114354 32274 115154
rect 34794 114354 34850 115154
rect 36726 114354 36782 115154
rect 38658 114354 38714 115154
rect 40590 114354 40646 115154
rect 43166 114354 43222 115154
rect 45098 114354 45154 115154
rect 47030 114354 47086 115154
rect 48962 114354 49018 115154
rect 51538 114354 51594 115154
rect 53470 114354 53526 115154
rect 55402 114354 55458 115154
rect 57334 114354 57390 115154
rect 59910 114354 59966 115154
rect 61842 114354 61898 115154
rect 63774 114354 63830 115154
rect 65706 114354 65762 115154
rect 68282 114354 68338 115154
rect 70214 114354 70270 115154
rect 72146 114354 72202 115154
rect 74078 114354 74134 115154
rect 76654 114354 76710 115154
rect 78586 114354 78642 115154
rect 80518 114354 80574 115154
rect 82450 114354 82506 115154
rect 85026 114354 85082 115154
rect 86958 114354 87014 115154
rect 88890 114354 88946 115154
rect 90822 114354 90878 115154
rect 93398 114354 93454 115154
rect 95330 114354 95386 115154
rect 97262 114354 97318 115154
rect 99194 114354 99250 115154
rect 101770 114354 101826 115154
rect 103702 114354 103758 115154
rect 105634 114354 105690 115154
rect 107566 114354 107622 115154
rect 110142 114354 110198 115154
rect 112074 114354 112130 115154
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 5814 0 5870 800
rect 7746 0 7802 800
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 14186 0 14242 800
rect 16118 0 16174 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 27066 0 27122 800
rect 28998 0 29054 800
rect 30930 0 30986 800
rect 32862 0 32918 800
rect 35438 0 35494 800
rect 37370 0 37426 800
rect 39302 0 39358 800
rect 41234 0 41290 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 49606 0 49662 800
rect 52182 0 52238 800
rect 54114 0 54170 800
rect 56046 0 56102 800
rect 57978 0 58034 800
rect 60554 0 60610 800
rect 62486 0 62542 800
rect 64418 0 64474 800
rect 66350 0 66406 800
rect 68926 0 68982 800
rect 70858 0 70914 800
rect 72790 0 72846 800
rect 74722 0 74778 800
rect 77298 0 77354 800
rect 79230 0 79286 800
rect 81162 0 81218 800
rect 83094 0 83150 800
rect 85670 0 85726 800
rect 87602 0 87658 800
rect 89534 0 89590 800
rect 91466 0 91522 800
rect 94042 0 94098 800
rect 95974 0 96030 800
rect 97906 0 97962 800
rect 99838 0 99894 800
rect 102414 0 102470 800
rect 104346 0 104402 800
rect 106278 0 106334 800
rect 108210 0 108266 800
rect 110786 0 110842 800
rect 112718 0 112774 800
<< obsm2 >>
rect 18 114298 1250 114458
rect 1418 114298 3182 114458
rect 3350 114298 5114 114458
rect 5282 114298 7046 114458
rect 7214 114298 9622 114458
rect 9790 114298 11554 114458
rect 11722 114298 13486 114458
rect 13654 114298 15418 114458
rect 15586 114298 17994 114458
rect 18162 114298 19926 114458
rect 20094 114298 21858 114458
rect 22026 114298 23790 114458
rect 23958 114298 26366 114458
rect 26534 114298 28298 114458
rect 28466 114298 30230 114458
rect 30398 114298 32162 114458
rect 32330 114298 34738 114458
rect 34906 114298 36670 114458
rect 36838 114298 38602 114458
rect 38770 114298 40534 114458
rect 40702 114298 43110 114458
rect 43278 114298 45042 114458
rect 45210 114298 46974 114458
rect 47142 114298 48906 114458
rect 49074 114298 51482 114458
rect 51650 114298 53414 114458
rect 53582 114298 55346 114458
rect 55514 114298 57278 114458
rect 57446 114298 59854 114458
rect 60022 114298 61786 114458
rect 61954 114298 63718 114458
rect 63886 114298 65650 114458
rect 65818 114298 68226 114458
rect 68394 114298 70158 114458
rect 70326 114298 72090 114458
rect 72258 114298 74022 114458
rect 74190 114298 76598 114458
rect 76766 114298 78530 114458
rect 78698 114298 80462 114458
rect 80630 114298 82394 114458
rect 82562 114298 84970 114458
rect 85138 114298 86902 114458
rect 87070 114298 88834 114458
rect 89002 114298 90766 114458
rect 90934 114298 93342 114458
rect 93510 114298 95274 114458
rect 95442 114298 97206 114458
rect 97374 114298 99138 114458
rect 99306 114298 101714 114458
rect 101882 114298 103646 114458
rect 103814 114298 105578 114458
rect 105746 114298 107510 114458
rect 107678 114298 110086 114458
rect 110254 114298 112018 114458
rect 112186 114298 112956 114458
rect 18 856 112956 114298
rect 130 734 1894 856
rect 2062 734 3826 856
rect 3994 734 5758 856
rect 5926 734 7690 856
rect 7858 734 10266 856
rect 10434 734 12198 856
rect 12366 734 14130 856
rect 14298 734 16062 856
rect 16230 734 18638 856
rect 18806 734 20570 856
rect 20738 734 22502 856
rect 22670 734 24434 856
rect 24602 734 27010 856
rect 27178 734 28942 856
rect 29110 734 30874 856
rect 31042 734 32806 856
rect 32974 734 35382 856
rect 35550 734 37314 856
rect 37482 734 39246 856
rect 39414 734 41178 856
rect 41346 734 43754 856
rect 43922 734 45686 856
rect 45854 734 47618 856
rect 47786 734 49550 856
rect 49718 734 52126 856
rect 52294 734 54058 856
rect 54226 734 55990 856
rect 56158 734 57922 856
rect 58090 734 60498 856
rect 60666 734 62430 856
rect 62598 734 64362 856
rect 64530 734 66294 856
rect 66462 734 68870 856
rect 69038 734 70802 856
rect 70970 734 72734 856
rect 72902 734 74666 856
rect 74834 734 77242 856
rect 77410 734 79174 856
rect 79342 734 81106 856
rect 81274 734 83038 856
rect 83206 734 85614 856
rect 85782 734 87546 856
rect 87714 734 89478 856
rect 89646 734 91410 856
rect 91578 734 93986 856
rect 94154 734 95918 856
rect 96086 734 97850 856
rect 98018 734 99782 856
rect 99950 734 102358 856
rect 102526 734 104290 856
rect 104458 734 106222 856
rect 106390 734 108154 856
rect 108322 734 110730 856
rect 110898 734 112662 856
rect 112830 734 112956 856
<< metal3 >>
rect 0 114248 800 114368
rect 112210 114248 113010 114368
rect 0 112208 800 112328
rect 112210 112208 113010 112328
rect 0 110168 800 110288
rect 112210 109488 113010 109608
rect 0 108128 800 108248
rect 112210 107448 113010 107568
rect 0 105408 800 105528
rect 112210 105408 113010 105528
rect 0 103368 800 103488
rect 112210 103368 113010 103488
rect 0 101328 800 101448
rect 112210 100648 113010 100768
rect 0 99288 800 99408
rect 112210 98608 113010 98728
rect 0 96568 800 96688
rect 112210 96568 113010 96688
rect 0 94528 800 94648
rect 112210 94528 113010 94648
rect 0 92488 800 92608
rect 112210 91808 113010 91928
rect 0 90448 800 90568
rect 112210 89768 113010 89888
rect 0 87728 800 87848
rect 112210 87728 113010 87848
rect 0 85688 800 85808
rect 112210 85688 113010 85808
rect 0 83648 800 83768
rect 112210 82968 113010 83088
rect 0 81608 800 81728
rect 112210 80928 113010 81048
rect 0 78888 800 79008
rect 112210 78888 113010 79008
rect 0 76848 800 76968
rect 112210 76848 113010 76968
rect 0 74808 800 74928
rect 112210 74128 113010 74248
rect 0 72768 800 72888
rect 112210 72088 113010 72208
rect 0 70048 800 70168
rect 112210 70048 113010 70168
rect 0 68008 800 68128
rect 112210 68008 113010 68128
rect 0 65968 800 66088
rect 112210 65288 113010 65408
rect 0 63928 800 64048
rect 112210 63248 113010 63368
rect 0 61208 800 61328
rect 112210 61208 113010 61328
rect 0 59168 800 59288
rect 112210 59168 113010 59288
rect 0 57128 800 57248
rect 112210 56448 113010 56568
rect 0 55088 800 55208
rect 112210 54408 113010 54528
rect 0 52368 800 52488
rect 112210 52368 113010 52488
rect 0 50328 800 50448
rect 112210 50328 113010 50448
rect 0 48288 800 48408
rect 112210 47608 113010 47728
rect 0 46248 800 46368
rect 112210 45568 113010 45688
rect 0 43528 800 43648
rect 112210 43528 113010 43648
rect 0 41488 800 41608
rect 112210 41488 113010 41608
rect 0 39448 800 39568
rect 112210 38768 113010 38888
rect 0 37408 800 37528
rect 112210 36728 113010 36848
rect 0 34688 800 34808
rect 112210 34688 113010 34808
rect 0 32648 800 32768
rect 112210 32648 113010 32768
rect 0 30608 800 30728
rect 112210 29928 113010 30048
rect 0 28568 800 28688
rect 112210 27888 113010 28008
rect 0 25848 800 25968
rect 112210 25848 113010 25968
rect 0 23808 800 23928
rect 112210 23808 113010 23928
rect 0 21768 800 21888
rect 112210 21088 113010 21208
rect 0 19728 800 19848
rect 112210 19048 113010 19168
rect 0 17008 800 17128
rect 112210 17008 113010 17128
rect 0 14968 800 15088
rect 112210 14968 113010 15088
rect 0 12928 800 13048
rect 112210 12248 113010 12368
rect 0 10888 800 11008
rect 112210 10208 113010 10328
rect 0 8168 800 8288
rect 112210 8168 113010 8288
rect 0 6128 800 6248
rect 112210 6128 113010 6248
rect 0 4088 800 4208
rect 112210 3408 113010 3528
rect 0 2048 800 2168
rect 112210 1368 113010 1488
<< obsm3 >>
rect 880 114168 112130 114341
rect 13 112408 112411 114168
rect 880 112128 112130 112408
rect 13 110368 112411 112128
rect 880 110088 112411 110368
rect 13 109688 112411 110088
rect 13 109408 112130 109688
rect 13 108328 112411 109408
rect 880 108048 112411 108328
rect 13 107648 112411 108048
rect 13 107368 112130 107648
rect 13 105608 112411 107368
rect 880 105328 112130 105608
rect 13 103568 112411 105328
rect 880 103288 112130 103568
rect 13 101528 112411 103288
rect 880 101248 112411 101528
rect 13 100848 112411 101248
rect 13 100568 112130 100848
rect 13 99488 112411 100568
rect 880 99208 112411 99488
rect 13 98808 112411 99208
rect 13 98528 112130 98808
rect 13 96768 112411 98528
rect 880 96488 112130 96768
rect 13 94728 112411 96488
rect 880 94448 112130 94728
rect 13 92688 112411 94448
rect 880 92408 112411 92688
rect 13 92008 112411 92408
rect 13 91728 112130 92008
rect 13 90648 112411 91728
rect 880 90368 112411 90648
rect 13 89968 112411 90368
rect 13 89688 112130 89968
rect 13 87928 112411 89688
rect 880 87648 112130 87928
rect 13 85888 112411 87648
rect 880 85608 112130 85888
rect 13 83848 112411 85608
rect 880 83568 112411 83848
rect 13 83168 112411 83568
rect 13 82888 112130 83168
rect 13 81808 112411 82888
rect 880 81528 112411 81808
rect 13 81128 112411 81528
rect 13 80848 112130 81128
rect 13 79088 112411 80848
rect 880 78808 112130 79088
rect 13 77048 112411 78808
rect 880 76768 112130 77048
rect 13 75008 112411 76768
rect 880 74728 112411 75008
rect 13 74328 112411 74728
rect 13 74048 112130 74328
rect 13 72968 112411 74048
rect 880 72688 112411 72968
rect 13 72288 112411 72688
rect 13 72008 112130 72288
rect 13 70248 112411 72008
rect 880 69968 112130 70248
rect 13 68208 112411 69968
rect 880 67928 112130 68208
rect 13 66168 112411 67928
rect 880 65888 112411 66168
rect 13 65488 112411 65888
rect 13 65208 112130 65488
rect 13 64128 112411 65208
rect 880 63848 112411 64128
rect 13 63448 112411 63848
rect 13 63168 112130 63448
rect 13 61408 112411 63168
rect 880 61128 112130 61408
rect 13 59368 112411 61128
rect 880 59088 112130 59368
rect 13 57328 112411 59088
rect 880 57048 112411 57328
rect 13 56648 112411 57048
rect 13 56368 112130 56648
rect 13 55288 112411 56368
rect 880 55008 112411 55288
rect 13 54608 112411 55008
rect 13 54328 112130 54608
rect 13 52568 112411 54328
rect 880 52288 112130 52568
rect 13 50528 112411 52288
rect 880 50248 112130 50528
rect 13 48488 112411 50248
rect 880 48208 112411 48488
rect 13 47808 112411 48208
rect 13 47528 112130 47808
rect 13 46448 112411 47528
rect 880 46168 112411 46448
rect 13 45768 112411 46168
rect 13 45488 112130 45768
rect 13 43728 112411 45488
rect 880 43448 112130 43728
rect 13 41688 112411 43448
rect 880 41408 112130 41688
rect 13 39648 112411 41408
rect 880 39368 112411 39648
rect 13 38968 112411 39368
rect 13 38688 112130 38968
rect 13 37608 112411 38688
rect 880 37328 112411 37608
rect 13 36928 112411 37328
rect 13 36648 112130 36928
rect 13 34888 112411 36648
rect 880 34608 112130 34888
rect 13 32848 112411 34608
rect 880 32568 112130 32848
rect 13 30808 112411 32568
rect 880 30528 112411 30808
rect 13 30128 112411 30528
rect 13 29848 112130 30128
rect 13 28768 112411 29848
rect 880 28488 112411 28768
rect 13 28088 112411 28488
rect 13 27808 112130 28088
rect 13 26048 112411 27808
rect 880 25768 112130 26048
rect 13 24008 112411 25768
rect 880 23728 112130 24008
rect 13 21968 112411 23728
rect 880 21688 112411 21968
rect 13 21288 112411 21688
rect 13 21008 112130 21288
rect 13 19928 112411 21008
rect 880 19648 112411 19928
rect 13 19248 112411 19648
rect 13 18968 112130 19248
rect 13 17208 112411 18968
rect 880 16928 112130 17208
rect 13 15168 112411 16928
rect 880 14888 112130 15168
rect 13 13128 112411 14888
rect 880 12848 112411 13128
rect 13 12448 112411 12848
rect 13 12168 112130 12448
rect 13 11088 112411 12168
rect 880 10808 112411 11088
rect 13 10408 112411 10808
rect 13 10128 112130 10408
rect 13 8368 112411 10128
rect 880 8088 112130 8368
rect 13 6328 112411 8088
rect 880 6048 112130 6328
rect 13 4288 112411 6048
rect 880 4008 112411 4288
rect 13 3608 112411 4008
rect 13 3328 112130 3608
rect 13 2248 112411 3328
rect 880 1968 112411 2248
rect 13 1568 112411 1968
rect 13 1395 112130 1568
<< metal4 >>
rect 4208 2128 4528 112656
rect 19568 2128 19888 112656
rect 34928 2128 35248 112656
rect 50288 2128 50608 112656
rect 65648 2128 65968 112656
rect 81008 2128 81328 112656
rect 96368 2128 96688 112656
<< obsm4 >>
rect 59 3299 4128 112437
rect 4608 3299 19488 112437
rect 19968 3299 34848 112437
rect 35328 3299 50208 112437
rect 50688 3299 65568 112437
rect 66048 3299 80928 112437
rect 81408 3299 96288 112437
rect 96768 3299 110893 112437
<< labels >>
rlabel metal2 s 37370 0 37426 800 6 active
port 1 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 112210 50328 113010 50448 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 112210 36728 113010 36848 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 26422 114354 26478 115154 6 io_in[15]
port 8 nsew signal input
rlabel metal3 s 112210 103368 113010 103488 6 io_in[16]
port 9 nsew signal input
rlabel metal3 s 112210 12248 113010 12368 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 13542 114354 13598 115154 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 97262 114354 97318 115154 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 19982 114354 20038 115154 6 io_in[24]
port 18 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 112210 34688 113010 34808 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 85026 114354 85082 115154 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 23846 114354 23902 115154 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 61842 114354 61898 115154 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 65706 114354 65762 115154 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 21914 114354 21970 115154 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 112210 98608 113010 98728 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 112210 68008 113010 68128 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 99194 114354 99250 115154 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 112074 114354 112130 115154 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 76654 114354 76710 115154 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 51538 114354 51594 115154 6 io_oeb[0]
port 40 nsew signal bidirectional
rlabel metal2 s 89534 0 89590 800 6 io_oeb[10]
port 41 nsew signal bidirectional
rlabel metal2 s 56046 0 56102 800 6 io_oeb[11]
port 42 nsew signal bidirectional
rlabel metal3 s 112210 72088 113010 72208 6 io_oeb[12]
port 43 nsew signal bidirectional
rlabel metal2 s 60554 0 60610 800 6 io_oeb[13]
port 44 nsew signal bidirectional
rlabel metal3 s 0 43528 800 43648 6 io_oeb[14]
port 45 nsew signal bidirectional
rlabel metal2 s 35438 0 35494 800 6 io_oeb[15]
port 46 nsew signal bidirectional
rlabel metal2 s 30286 114354 30342 115154 6 io_oeb[16]
port 47 nsew signal bidirectional
rlabel metal3 s 112210 8168 113010 8288 6 io_oeb[17]
port 48 nsew signal bidirectional
rlabel metal2 s 15474 114354 15530 115154 6 io_oeb[18]
port 49 nsew signal bidirectional
rlabel metal3 s 0 17008 800 17128 6 io_oeb[19]
port 50 nsew signal bidirectional
rlabel metal3 s 112210 74128 113010 74248 6 io_oeb[1]
port 51 nsew signal bidirectional
rlabel metal2 s 91466 0 91522 800 6 io_oeb[20]
port 52 nsew signal bidirectional
rlabel metal3 s 112210 109488 113010 109608 6 io_oeb[21]
port 53 nsew signal bidirectional
rlabel metal3 s 0 70048 800 70168 6 io_oeb[22]
port 54 nsew signal bidirectional
rlabel metal2 s 12254 0 12310 800 6 io_oeb[23]
port 55 nsew signal bidirectional
rlabel metal2 s 55402 114354 55458 115154 6 io_oeb[24]
port 56 nsew signal bidirectional
rlabel metal3 s 112210 32648 113010 32768 6 io_oeb[25]
port 57 nsew signal bidirectional
rlabel metal2 s 110786 0 110842 800 6 io_oeb[26]
port 58 nsew signal bidirectional
rlabel metal3 s 112210 91808 113010 91928 6 io_oeb[27]
port 59 nsew signal bidirectional
rlabel metal3 s 112210 114248 113010 114368 6 io_oeb[28]
port 60 nsew signal bidirectional
rlabel metal2 s 97906 0 97962 800 6 io_oeb[29]
port 61 nsew signal bidirectional
rlabel metal3 s 112210 76848 113010 76968 6 io_oeb[2]
port 62 nsew signal bidirectional
rlabel metal3 s 112210 52368 113010 52488 6 io_oeb[30]
port 63 nsew signal bidirectional
rlabel metal2 s 63774 114354 63830 115154 6 io_oeb[31]
port 64 nsew signal bidirectional
rlabel metal3 s 112210 61208 113010 61328 6 io_oeb[32]
port 65 nsew signal bidirectional
rlabel metal3 s 0 41488 800 41608 6 io_oeb[33]
port 66 nsew signal bidirectional
rlabel metal2 s 40590 114354 40646 115154 6 io_oeb[34]
port 67 nsew signal bidirectional
rlabel metal2 s 57334 114354 57390 115154 6 io_oeb[35]
port 68 nsew signal bidirectional
rlabel metal3 s 0 50328 800 50448 6 io_oeb[36]
port 69 nsew signal bidirectional
rlabel metal3 s 0 25848 800 25968 6 io_oeb[37]
port 70 nsew signal bidirectional
rlabel metal3 s 0 101328 800 101448 6 io_oeb[3]
port 71 nsew signal bidirectional
rlabel metal3 s 0 39448 800 39568 6 io_oeb[4]
port 72 nsew signal bidirectional
rlabel metal3 s 112210 3408 113010 3528 6 io_oeb[5]
port 73 nsew signal bidirectional
rlabel metal3 s 0 74808 800 74928 6 io_oeb[6]
port 74 nsew signal bidirectional
rlabel metal3 s 112210 43528 113010 43648 6 io_oeb[7]
port 75 nsew signal bidirectional
rlabel metal2 s 28354 114354 28410 115154 6 io_oeb[8]
port 76 nsew signal bidirectional
rlabel metal2 s 10322 0 10378 800 6 io_oeb[9]
port 77 nsew signal bidirectional
rlabel metal2 s 24490 0 24546 800 6 io_out[0]
port 78 nsew signal bidirectional
rlabel metal2 s 93398 114354 93454 115154 6 io_out[10]
port 79 nsew signal bidirectional
rlabel metal3 s 112210 65288 113010 65408 6 io_out[11]
port 80 nsew signal bidirectional
rlabel metal3 s 0 6128 800 6248 6 io_out[12]
port 81 nsew signal bidirectional
rlabel metal3 s 0 14968 800 15088 6 io_out[13]
port 82 nsew signal bidirectional
rlabel metal2 s 94042 0 94098 800 6 io_out[14]
port 83 nsew signal bidirectional
rlabel metal3 s 0 85688 800 85808 6 io_out[15]
port 84 nsew signal bidirectional
rlabel metal3 s 0 94528 800 94648 6 io_out[16]
port 85 nsew signal bidirectional
rlabel metal3 s 112210 63248 113010 63368 6 io_out[17]
port 86 nsew signal bidirectional
rlabel metal2 s 32218 114354 32274 115154 6 io_out[18]
port 87 nsew signal bidirectional
rlabel metal3 s 112210 94528 113010 94648 6 io_out[19]
port 88 nsew signal bidirectional
rlabel metal3 s 112210 41488 113010 41608 6 io_out[1]
port 89 nsew signal bidirectional
rlabel metal2 s 99838 0 99894 800 6 io_out[20]
port 90 nsew signal bidirectional
rlabel metal2 s 90822 114354 90878 115154 6 io_out[21]
port 91 nsew signal bidirectional
rlabel metal3 s 0 92488 800 92608 6 io_out[22]
port 92 nsew signal bidirectional
rlabel metal2 s 74722 0 74778 800 6 io_out[23]
port 93 nsew signal bidirectional
rlabel metal3 s 0 2048 800 2168 6 io_out[24]
port 94 nsew signal bidirectional
rlabel metal2 s 62486 0 62542 800 6 io_out[25]
port 95 nsew signal bidirectional
rlabel metal2 s 82450 114354 82506 115154 6 io_out[26]
port 96 nsew signal bidirectional
rlabel metal2 s 68282 114354 68338 115154 6 io_out[27]
port 97 nsew signal bidirectional
rlabel metal2 s 86958 114354 87014 115154 6 io_out[28]
port 98 nsew signal bidirectional
rlabel metal2 s 39302 0 39358 800 6 io_out[29]
port 99 nsew signal bidirectional
rlabel metal3 s 112210 6128 113010 6248 6 io_out[2]
port 100 nsew signal bidirectional
rlabel metal2 s 16118 0 16174 800 6 io_out[30]
port 101 nsew signal bidirectional
rlabel metal3 s 0 65968 800 66088 6 io_out[31]
port 102 nsew signal bidirectional
rlabel metal2 s 103702 114354 103758 115154 6 io_out[32]
port 103 nsew signal bidirectional
rlabel metal3 s 0 108128 800 108248 6 io_out[33]
port 104 nsew signal bidirectional
rlabel metal3 s 112210 17008 113010 17128 6 io_out[34]
port 105 nsew signal bidirectional
rlabel metal3 s 112210 96568 113010 96688 6 io_out[35]
port 106 nsew signal bidirectional
rlabel metal3 s 112210 89768 113010 89888 6 io_out[36]
port 107 nsew signal bidirectional
rlabel metal2 s 34794 114354 34850 115154 6 io_out[37]
port 108 nsew signal bidirectional
rlabel metal3 s 112210 105408 113010 105528 6 io_out[3]
port 109 nsew signal bidirectional
rlabel metal2 s 74078 114354 74134 115154 6 io_out[4]
port 110 nsew signal bidirectional
rlabel metal3 s 112210 70048 113010 70168 6 io_out[5]
port 111 nsew signal bidirectional
rlabel metal3 s 112210 87728 113010 87848 6 io_out[6]
port 112 nsew signal bidirectional
rlabel metal2 s 107566 114354 107622 115154 6 io_out[7]
port 113 nsew signal bidirectional
rlabel metal3 s 0 46248 800 46368 6 io_out[8]
port 114 nsew signal bidirectional
rlabel metal2 s 43810 0 43866 800 6 io_out[9]
port 115 nsew signal bidirectional
rlabel metal3 s 112210 23808 113010 23928 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal3 s 112210 19048 113010 19168 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal2 s 3238 114354 3294 115154 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 36726 114354 36782 115154 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 53470 114354 53526 115154 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 38658 114354 38714 115154 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal2 s 110142 114354 110198 115154 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal3 s 112210 21088 113010 21208 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal3 s 112210 56448 113010 56568 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 112210 10208 113010 10328 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal2 s 1306 114354 1362 115154 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal2 s 9678 114354 9734 115154 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal2 s 95330 114354 95386 115154 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 5170 114354 5226 115154 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal2 s 43166 114354 43222 115154 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal2 s 45098 114354 45154 115154 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 la1_data_out[0]
port 148 nsew signal bidirectional
rlabel metal2 s 18694 0 18750 800 6 la1_data_out[10]
port 149 nsew signal bidirectional
rlabel metal3 s 112210 27888 113010 28008 6 la1_data_out[11]
port 150 nsew signal bidirectional
rlabel metal2 s 52182 0 52238 800 6 la1_data_out[12]
port 151 nsew signal bidirectional
rlabel metal3 s 112210 107448 113010 107568 6 la1_data_out[13]
port 152 nsew signal bidirectional
rlabel metal3 s 112210 82968 113010 83088 6 la1_data_out[14]
port 153 nsew signal bidirectional
rlabel metal2 s 59910 114354 59966 115154 6 la1_data_out[15]
port 154 nsew signal bidirectional
rlabel metal3 s 0 96568 800 96688 6 la1_data_out[16]
port 155 nsew signal bidirectional
rlabel metal3 s 112210 38768 113010 38888 6 la1_data_out[17]
port 156 nsew signal bidirectional
rlabel metal3 s 0 76848 800 76968 6 la1_data_out[18]
port 157 nsew signal bidirectional
rlabel metal2 s 11610 114354 11666 115154 6 la1_data_out[19]
port 158 nsew signal bidirectional
rlabel metal3 s 112210 59168 113010 59288 6 la1_data_out[1]
port 159 nsew signal bidirectional
rlabel metal3 s 0 103368 800 103488 6 la1_data_out[20]
port 160 nsew signal bidirectional
rlabel metal2 s 66350 0 66406 800 6 la1_data_out[21]
port 161 nsew signal bidirectional
rlabel metal3 s 112210 100648 113010 100768 6 la1_data_out[22]
port 162 nsew signal bidirectional
rlabel metal2 s 70214 114354 70270 115154 6 la1_data_out[23]
port 163 nsew signal bidirectional
rlabel metal2 s 28998 0 29054 800 6 la1_data_out[24]
port 164 nsew signal bidirectional
rlabel metal3 s 112210 45568 113010 45688 6 la1_data_out[25]
port 165 nsew signal bidirectional
rlabel metal3 s 0 8168 800 8288 6 la1_data_out[26]
port 166 nsew signal bidirectional
rlabel metal3 s 112210 14968 113010 15088 6 la1_data_out[27]
port 167 nsew signal bidirectional
rlabel metal3 s 0 110168 800 110288 6 la1_data_out[28]
port 168 nsew signal bidirectional
rlabel metal2 s 102414 0 102470 800 6 la1_data_out[29]
port 169 nsew signal bidirectional
rlabel metal2 s 14186 0 14242 800 6 la1_data_out[2]
port 170 nsew signal bidirectional
rlabel metal2 s 47674 0 47730 800 6 la1_data_out[30]
port 171 nsew signal bidirectional
rlabel metal3 s 112210 29928 113010 30048 6 la1_data_out[31]
port 172 nsew signal bidirectional
rlabel metal3 s 112210 112208 113010 112328 6 la1_data_out[3]
port 173 nsew signal bidirectional
rlabel metal3 s 0 30608 800 30728 6 la1_data_out[4]
port 174 nsew signal bidirectional
rlabel metal2 s 104346 0 104402 800 6 la1_data_out[5]
port 175 nsew signal bidirectional
rlabel metal2 s 7746 0 7802 800 6 la1_data_out[6]
port 176 nsew signal bidirectional
rlabel metal3 s 112210 47608 113010 47728 6 la1_data_out[7]
port 177 nsew signal bidirectional
rlabel metal2 s 1950 0 2006 800 6 la1_data_out[8]
port 178 nsew signal bidirectional
rlabel metal3 s 112210 85688 113010 85808 6 la1_data_out[9]
port 179 nsew signal bidirectional
rlabel metal2 s 105634 114354 105690 115154 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 112210 1368 113010 1488 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal2 s 101770 114354 101826 115154 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal2 s 18 0 74 800 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal2 s 7102 114354 7158 115154 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal2 s 48962 114354 49018 115154 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal2 s 72146 114354 72202 115154 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal2 s 47030 114354 47086 115154 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal2 s 88890 114354 88946 115154 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 112210 25848 113010 25968 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 112210 80928 113010 81048 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 112210 78888 113010 79008 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal2 s 80518 114354 80574 115154 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal2 s 78586 114354 78642 115154 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal2 s 18050 114354 18106 115154 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 user_clock2
port 212 nsew signal input
rlabel metal4 s 4208 2128 4528 112656 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 112656 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 112656 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 112656 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 112656 6 vssd1
port 214 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 112656 6 vssd1
port 214 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 112656 6 vssd1
port 214 nsew ground bidirectional
rlabel metal3 s 112210 54408 113010 54528 6 wb_clk_i
port 215 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 113010 115154
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 49101584
string GDS_FILE /openlane/designs/wrapped_ibnalhaytham/runs/RUN_2022.08.27_14.16.49/results/signoff/wrapped_ibnalhaytham.magic.gds
string GDS_START 966832
<< end >>

